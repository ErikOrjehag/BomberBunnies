library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_000111100101", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000110010100", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011000100", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000010000", -- BOOM1
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000001101010", -- BOOM2
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  16 => b"00000_0000_00_001010000111", -- load, gr0, P1EXPLOSION1ACTIVE
  17 => b"00011_0000_01_000000000000", -- sub, gr0
  18 => b"00000_0000_00_000000000001", -- 1
  19 => b"00111_0000_01_000000000000", -- bne
  20 => b"00000_0000_00_000000001100", -- BOOM1_R
  21 => b"00000_0000_00_001010000110", -- load, gr0, P1EXPLOSION1TIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000001", -- 1
  24 => b"00001_0000_10_001010000110", -- store, gr0, P1EXPLOSION1TIME
  25 => b"00000_0000_00_001010000110", -- load, gr0, P1EXPLOSION1TIME
  26 => b"00011_0000_01_000000000000", -- sub, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00111_0000_01_000000000000", -- bne
  29 => b"00000_0000_00_000000001100", -- BOOM1_R
  30 => b"00000_0000_01_000000000000", -- load, gr0
  31 => b"00000_0000_00_000000000000", -- 0
  32 => b"00001_0000_10_001010000111", -- store, gr0, P1EXPLOSION1ACTIVE
  33 => b"00000_0010_00_001010001000", -- load, gr2, P1EXPLOSION1POS
  34 => b"00000_0011_00_001010110001", -- load, gr3, GRASS
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01110_0011_00_000000000000", -- twrite, gr3
  37 => b"00010_0010_01_000000000000", -- add, gr2
  38 => b"00000_0000_00_000000000001", -- 1
  39 => b"10000_0010_00_000000000000", -- tpoint, gr2
  40 => b"01111_0000_00_000000000000", -- tread, gr0
  41 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  42 => b"00111_0000_01_000000000000", -- bne
  43 => b"00000_0000_00_000000110101", -- E1LEFT
  44 => b"01110_0011_00_000000000000", -- twrite, gr3
  45 => b"00010_0010_01_000000000000", -- add, gr2
  46 => b"00000_0000_00_000000000001", -- 1
  47 => b"10000_0010_00_000000000000", -- tpoint, gr2
  48 => b"01111_0000_00_000000000000", -- tread, gr0
  49 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  50 => b"00111_0000_01_000000000000", -- bne
  51 => b"00000_0000_00_000000110101", -- E1LEFT
  52 => b"01110_0011_00_000000000000", -- twrite, gr3
  53 => b"00000_0010_00_001010001000", -- load, gr2, P1EXPLOSION1POS
  54 => b"00011_0010_01_000000000000", -- sub, gr2
  55 => b"00000_0000_00_000000000001", -- 1
  56 => b"10000_0010_00_000000000000", -- tpoint, gr2
  57 => b"01111_0000_00_000000000000", -- tread, gr0
  58 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  59 => b"00111_0000_01_000000000000", -- bne
  60 => b"00000_0000_00_000001000110", -- E1DOWN
  61 => b"01110_0011_00_000000000000", -- twrite, gr3
  62 => b"00011_0010_01_000000000000", -- sub, gr2
  63 => b"00000_0000_00_000000000001", -- 1
  64 => b"10000_0010_00_000000000000", -- tpoint, gr2
  65 => b"01111_0000_00_000000000000", -- tread, gr0
  66 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  67 => b"00111_0000_01_000000000000", -- bne
  68 => b"00000_0000_00_000001000110", -- E1DOWN
  69 => b"01110_0011_00_000000000000", -- twrite, gr3
  70 => b"00000_0010_00_001010001000", -- load, gr2, P1EXPLOSION1POS
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000001111", -- 15
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0000_00_000000000000", -- tread, gr0
  75 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  76 => b"00111_0000_01_000000000000", -- bne
  77 => b"00000_0000_00_000001010111", -- E1UP
  78 => b"01110_0011_00_000000000000", -- twrite, gr3
  79 => b"00010_0010_01_000000000000", -- add, gr2
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"10000_0010_00_000000000000", -- tpoint, gr2
  82 => b"01111_0000_00_000000000000", -- tread, gr0
  83 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  84 => b"00111_0000_01_000000000000", -- bne
  85 => b"00000_0000_00_000001010111", -- E1UP
  86 => b"01110_0011_00_000000000000", -- twrite, gr3
  87 => b"00000_0010_00_001010001000", -- load, gr2, P1EXPLOSION1POS
  88 => b"00011_0010_01_000000000000", -- sub, gr2
  89 => b"00000_0000_00_000000001111", -- 15
  90 => b"10000_0010_00_000000000000", -- tpoint, gr2
  91 => b"01111_0000_00_000000000000", -- tread, gr0
  92 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
  93 => b"00111_0000_01_000000000000", -- bne
  94 => b"00000_0000_00_000000001100", -- BOOM1_R
  95 => b"01110_0011_00_000000000000", -- twrite, gr3
  96 => b"00011_0010_01_000000000000", -- sub, gr2
  97 => b"00000_0000_00_000000001111", -- 15
  98 => b"10000_0010_00_000000000000", -- tpoint, gr2
  99 => b"01111_0000_00_000000000000", -- tread, gr0
 100 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 101 => b"00111_0000_01_000000000000", -- bne
 102 => b"00000_0000_00_000000001100", -- BOOM1_R
 103 => b"01110_0011_00_000000000000", -- twrite, gr3
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000000001100", -- BOOM1_R
 106 => b"00000_0000_00_001010011001", -- load, gr0, P2EXPLOSION4ACTIVE
 107 => b"00011_0000_01_000000000000", -- sub, gr0
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00111_0000_01_000000000000", -- bne
 110 => b"00000_0000_00_000000001110", -- BOOM2_R
 111 => b"00000_0000_00_001010011000", -- load, gr0, P2EXPLOSION4TIME
 112 => b"00011_0000_01_000000000000", -- sub, gr0
 113 => b"00000_0000_00_000000000001", -- 1
 114 => b"00001_0000_10_001010011000", -- store, gr0, P2EXPLOSION4TIME
 115 => b"00000_0000_00_001010011000", -- load, gr0, P2EXPLOSION4TIME
 116 => b"00011_0000_01_000000000000", -- sub, gr0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00111_0000_01_000000000000", -- bne
 119 => b"00000_0000_00_000000001110", -- BOOM2_R
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001010011001", -- store, gr0, P2EXPLOSION4ACTIVE
 123 => b"00000_0010_00_001010011010", -- load, gr2, P2EXPLOSION4POS
 124 => b"00000_0011_00_001010110001", -- load, gr3, GRASS
 125 => b"10000_0010_00_000000000000", -- tpoint, gr2
 126 => b"01110_0011_00_000000000000", -- twrite, gr3
 127 => b"00010_0010_01_000000000000", -- add, gr2
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"10000_0010_00_000000000000", -- tpoint, gr2
 130 => b"01111_0000_00_000000000000", -- tread, gr0
 131 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 132 => b"00111_0000_01_000000000000", -- bne
 133 => b"00000_0000_00_000010001111", -- E2LEFT
 134 => b"01110_0011_00_000000000000", -- twrite, gr3
 135 => b"00010_0010_01_000000000000", -- add, gr2
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0010_00_000000000000", -- tpoint, gr2
 138 => b"01111_0000_00_000000000000", -- tread, gr0
 139 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000010001111", -- E2LEFT
 142 => b"01110_0011_00_000000000000", -- twrite, gr3
 143 => b"00000_0010_00_001010011010", -- load, gr2, P2EXPLOSION4POS
 144 => b"00011_0010_01_000000000000", -- sub, gr2
 145 => b"00000_0000_00_000000000001", -- 1
 146 => b"10000_0010_00_000000000000", -- tpoint, gr2
 147 => b"01111_0000_00_000000000000", -- tread, gr0
 148 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 149 => b"00111_0000_01_000000000000", -- bne
 150 => b"00000_0000_00_000010100000", -- E2DOWN
 151 => b"01110_0011_00_000000000000", -- twrite, gr3
 152 => b"00011_0010_01_000000000000", -- sub, gr2
 153 => b"00000_0000_00_000000000001", -- 1
 154 => b"10000_0010_00_000000000000", -- tpoint, gr2
 155 => b"01111_0000_00_000000000000", -- tread, gr0
 156 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000010100000", -- E2DOWN
 159 => b"01110_0011_00_000000000000", -- twrite, gr3
 160 => b"00000_0010_00_001010011010", -- load, gr2, P2EXPLOSION4POS
 161 => b"00010_0010_01_000000000000", -- add, gr2
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"10000_0010_00_000000000000", -- tpoint, gr2
 164 => b"01111_0000_00_000000000000", -- tread, gr0
 165 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 166 => b"00111_0000_01_000000000000", -- bne
 167 => b"00000_0000_00_000010110001", -- E2UP
 168 => b"01110_0011_00_000000000000", -- twrite, gr3
 169 => b"00010_0010_01_000000000000", -- add, gr2
 170 => b"00000_0000_00_000000001111", -- 15
 171 => b"10000_0010_00_000000000000", -- tpoint, gr2
 172 => b"01111_0000_00_000000000000", -- tread, gr0
 173 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000010110001", -- E2UP
 176 => b"01110_0011_00_000000000000", -- twrite, gr3
 177 => b"00000_0010_00_001010011010", -- load, gr2, P2EXPLOSION4POS
 178 => b"00011_0010_01_000000000000", -- sub, gr2
 179 => b"00000_0000_00_000000001111", -- 15
 180 => b"10000_0010_00_000000000000", -- tpoint, gr2
 181 => b"01111_0000_00_000000000000", -- tread, gr0
 182 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 183 => b"00111_0000_01_000000000000", -- bne
 184 => b"00000_0000_00_000000001110", -- BOOM2_R
 185 => b"01110_0011_00_000000000000", -- twrite, gr3
 186 => b"00011_0010_01_000000000000", -- sub, gr2
 187 => b"00000_0000_00_000000001111", -- 15
 188 => b"10000_0010_00_000000000000", -- tpoint, gr2
 189 => b"01111_0000_00_000000000000", -- tread, gr0
 190 => b"00011_0000_00_001010110100", -- sub, gr0, EXPLOSION
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000001110", -- BOOM2_R
 193 => b"01110_0011_00_000000000000", -- twrite, gr3
 194 => b"00100_0000_01_000000000000", -- jump
 195 => b"00000_0000_00_000000001110", -- BOOM2_R
 196 => b"00100_0000_01_000000000000", -- jump
 197 => b"00000_0000_00_000011001010", -- TICKBOMB1
 198 => b"00100_0000_01_000000000000", -- jump
 199 => b"00000_0000_00_000100101111", -- TICKBOMB2
 200 => b"00100_0000_01_000000000000", -- jump
 201 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 202 => b"00000_0000_00_001010000101", -- load, gr0, P1BOMB1ACTIVE
 203 => b"00011_0000_01_000000000000", -- sub, gr0
 204 => b"00000_0000_00_000000000001", -- 1
 205 => b"00111_0000_01_000000000000", -- bne
 206 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 207 => b"00000_0000_00_001010000100", -- load, gr0, P1BOMB1TIME
 208 => b"00011_0000_01_000000000000", -- sub, gr0
 209 => b"00000_0000_00_000000000001", -- 1
 210 => b"00001_0000_10_001010000100", -- store, gr0, P1BOMB1TIME
 211 => b"00000_0000_01_000000000000", -- load, gr0
 212 => b"00000_0000_00_000000000000", -- 0
 213 => b"00011_0000_00_001010000100", -- sub, gr0, P1BOMB1TIME
 214 => b"00110_0000_01_000000000000", -- beq
 215 => b"00000_0000_00_000011011010", -- EXPLODE1
 216 => b"00100_0000_01_000000000000", -- jump
 217 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 218 => b"00000_0000_00_001010000011", -- load, gr0, P1BOMB1POS
 219 => b"00001_0000_10_001010001000", -- store, gr0, P1EXPLOSION1POS
 220 => b"00000_0000_01_000000000000", -- load, gr0
 221 => b"00000_0000_00_000000000001", -- 1
 222 => b"00001_0000_10_001010000111", -- store, gr0, P1EXPLOSION1ACTIVE
 223 => b"00000_0000_01_000000000000", -- load, gr0
 224 => b"00000_0000_00_000000000010", -- 2
 225 => b"00001_0000_10_001010000110", -- store, gr0, P1EXPLOSION1TIME
 226 => b"00000_0000_00_001010100111", -- load, gr0, P1BOMBCOUNT
 227 => b"00011_0000_01_000000000000", -- sub, gr0
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00001_0000_10_001010100111", -- store, gr0, P1BOMBCOUNT
 230 => b"00000_0010_00_001010000011", -- load, gr2, P1BOMB1POS
 231 => b"00000_0011_00_001010110100", -- load, gr3, EXPLOSION
 232 => b"10000_0010_00_000000000000", -- tpoint, gr2
 233 => b"01110_0011_00_000000000000", -- twrite, gr3
 234 => b"00010_0010_01_000000000000", -- add, gr2
 235 => b"00000_0000_00_000000000001", -- 1
 236 => b"10000_0010_00_000000000000", -- tpoint, gr2
 237 => b"01111_0000_00_000000000000", -- tread, gr0
 238 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 239 => b"00110_0000_01_000000000000", -- beq
 240 => b"00000_0000_00_000011111010", -- P1LEFT
 241 => b"01110_0011_00_000000000000", -- twrite, gr3
 242 => b"00010_0010_01_000000000000", -- add, gr2
 243 => b"00000_0000_00_000000000001", -- 1
 244 => b"10000_0010_00_000000000000", -- tpoint, gr2
 245 => b"01111_0000_00_000000000000", -- tread, gr0
 246 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 247 => b"00110_0000_01_000000000000", -- beq
 248 => b"00000_0000_00_000011111010", -- P1LEFT
 249 => b"01110_0011_00_000000000000", -- twrite, gr3
 250 => b"00000_0010_00_001010000011", -- load, gr2, P1BOMB1POS
 251 => b"00011_0010_01_000000000000", -- sub, gr2
 252 => b"00000_0000_00_000000000001", -- 1
 253 => b"10000_0010_00_000000000000", -- tpoint, gr2
 254 => b"01111_0000_00_000000000000", -- tread, gr0
 255 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 256 => b"00110_0000_01_000000000000", -- beq
 257 => b"00000_0000_00_000100001011", -- P1DOWN
 258 => b"01110_0011_00_000000000000", -- twrite, gr3
 259 => b"00011_0010_01_000000000000", -- sub, gr2
 260 => b"00000_0000_00_000000000001", -- 1
 261 => b"10000_0010_00_000000000000", -- tpoint, gr2
 262 => b"01111_0000_00_000000000000", -- tread, gr0
 263 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 264 => b"00110_0000_01_000000000000", -- beq
 265 => b"00000_0000_00_000100001011", -- P1DOWN
 266 => b"01110_0011_00_000000000000", -- twrite, gr3
 267 => b"00000_0010_00_001010000011", -- load, gr2, P1BOMB1POS
 268 => b"00010_0010_01_000000000000", -- add, gr2
 269 => b"00000_0000_00_000000001111", -- 15
 270 => b"10000_0010_00_000000000000", -- tpoint, gr2
 271 => b"01111_0000_00_000000000000", -- tread, gr0
 272 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 273 => b"00110_0000_01_000000000000", -- beq
 274 => b"00000_0000_00_000100011100", -- P1UP
 275 => b"01110_0011_00_000000000000", -- twrite, gr3
 276 => b"00010_0010_01_000000000000", -- add, gr2
 277 => b"00000_0000_00_000000001111", -- 15
 278 => b"10000_0010_00_000000000000", -- tpoint, gr2
 279 => b"01111_0000_00_000000000000", -- tread, gr0
 280 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 281 => b"00110_0000_01_000000000000", -- beq
 282 => b"00000_0000_00_000100011100", -- P1UP
 283 => b"01110_0011_00_000000000000", -- twrite, gr3
 284 => b"00000_0010_00_001010000011", -- load, gr2, P1BOMB1POS
 285 => b"00011_0010_01_000000000000", -- sub, gr2
 286 => b"00000_0000_00_000000001111", -- 15
 287 => b"10000_0010_00_000000000000", -- tpoint, gr2
 288 => b"01111_0000_00_000000000000", -- tread, gr0
 289 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 290 => b"00110_0000_01_000000000000", -- beq
 291 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 292 => b"01110_0011_00_000000000000", -- twrite, gr3
 293 => b"00011_0010_01_000000000000", -- sub, gr2
 294 => b"00000_0000_00_000000001111", -- 15
 295 => b"10000_0010_00_000000000000", -- tpoint, gr2
 296 => b"01111_0000_00_000000000000", -- tread, gr0
 297 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 298 => b"00110_0000_01_000000000000", -- beq
 299 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 300 => b"01110_0011_00_000000000000", -- twrite, gr3
 301 => b"00100_0000_01_000000000000", -- jump
 302 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 303 => b"00000_0000_00_001010010111", -- load, gr0, P2BOMB4ACTIVE
 304 => b"00011_0000_01_000000000000", -- sub, gr0
 305 => b"00000_0000_00_000000000001", -- 1
 306 => b"00111_0000_01_000000000000", -- bne
 307 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 308 => b"00000_0000_00_001010010110", -- load, gr0, P2BOMB4TIME
 309 => b"00011_0000_01_000000000000", -- sub, gr0
 310 => b"00000_0000_00_000000000001", -- 1
 311 => b"00001_0000_10_001010010110", -- store, gr0, P2BOMB4TIME
 312 => b"00000_0000_01_000000000000", -- load, gr0
 313 => b"00000_0000_00_000000000000", -- 0
 314 => b"00011_0000_00_001010010110", -- sub, gr0, P2BOMB4TIME
 315 => b"00110_0000_01_000000000000", -- beq
 316 => b"00000_0000_00_000100111111", -- EXPLODE2
 317 => b"00100_0000_01_000000000000", -- jump
 318 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 319 => b"00000_0000_00_001010010101", -- load, gr0, P2BOMB4POS
 320 => b"00001_0000_10_001010011010", -- store, gr0, P2EXPLOSION4POS
 321 => b"00000_0000_01_000000000000", -- load, gr0
 322 => b"00000_0000_00_000000000001", -- 1
 323 => b"00001_0000_10_001010011001", -- store, gr0, P2EXPLOSION4ACTIVE
 324 => b"00000_0000_01_000000000000", -- load, gr0
 325 => b"00000_0000_00_000000000010", -- 2
 326 => b"00001_0000_10_001010011000", -- store, gr0, P2EXPLOSION4TIME
 327 => b"00000_0000_00_001010101000", -- load, gr0, P2BOMBCOUNT
 328 => b"00011_0000_01_000000000000", -- sub, gr0
 329 => b"00000_0000_00_000000000001", -- 1
 330 => b"00001_0000_10_001010101000", -- store, gr0, P2BOMBCOUNT
 331 => b"00000_0010_00_001010010101", -- load, gr2, P2BOMB4POS
 332 => b"00000_0011_00_001010110100", -- load, gr3, EXPLOSION
 333 => b"10000_0010_00_000000000000", -- tpoint, gr2
 334 => b"01110_0011_00_000000000000", -- twrite, gr3
 335 => b"00010_0010_01_000000000000", -- add, gr2
 336 => b"00000_0000_00_000000000001", -- 1
 337 => b"10000_0010_00_000000000000", -- tpoint, gr2
 338 => b"01111_0000_00_000000000000", -- tread, gr0
 339 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 340 => b"00110_0000_01_000000000000", -- beq
 341 => b"00000_0000_00_000101011111", -- P2LEFT
 342 => b"01110_0011_00_000000000000", -- twrite, gr3
 343 => b"00010_0010_01_000000000000", -- add, gr2
 344 => b"00000_0000_00_000000000001", -- 1
 345 => b"10000_0010_00_000000000000", -- tpoint, gr2
 346 => b"01111_0000_00_000000000000", -- tread, gr0
 347 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 348 => b"00110_0000_01_000000000000", -- beq
 349 => b"00000_0000_00_000101011111", -- P2LEFT
 350 => b"01110_0011_00_000000000000", -- twrite, gr3
 351 => b"00000_0010_00_001010010101", -- load, gr2, P2BOMB4POS
 352 => b"00011_0010_01_000000000000", -- sub, gr2
 353 => b"00000_0000_00_000000000001", -- 1
 354 => b"10000_0010_00_000000000000", -- tpoint, gr2
 355 => b"01111_0000_00_000000000000", -- tread, gr0
 356 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 357 => b"00110_0000_01_000000000000", -- beq
 358 => b"00000_0000_00_000101110000", -- P2DOWN
 359 => b"01110_0011_00_000000000000", -- twrite, gr3
 360 => b"00011_0010_01_000000000000", -- sub, gr2
 361 => b"00000_0000_00_000000000001", -- 1
 362 => b"10000_0010_00_000000000000", -- tpoint, gr2
 363 => b"01111_0000_00_000000000000", -- tread, gr0
 364 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 365 => b"00110_0000_01_000000000000", -- beq
 366 => b"00000_0000_00_000101110000", -- P2DOWN
 367 => b"01110_0011_00_000000000000", -- twrite, gr3
 368 => b"00000_0010_00_001010010101", -- load, gr2, P2BOMB4POS
 369 => b"00010_0010_01_000000000000", -- add, gr2
 370 => b"00000_0000_00_000000001111", -- 15
 371 => b"10000_0010_00_000000000000", -- tpoint, gr2
 372 => b"01111_0000_00_000000000000", -- tread, gr0
 373 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 374 => b"00110_0000_01_000000000000", -- beq
 375 => b"00000_0000_00_000110000001", -- P2UP
 376 => b"01110_0011_00_000000000000", -- twrite, gr3
 377 => b"00010_0010_01_000000000000", -- add, gr2
 378 => b"00000_0000_00_000000001111", -- 15
 379 => b"10000_0010_00_000000000000", -- tpoint, gr2
 380 => b"01111_0000_00_000000000000", -- tread, gr0
 381 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 382 => b"00110_0000_01_000000000000", -- beq
 383 => b"00000_0000_00_000110000001", -- P2UP
 384 => b"01110_0011_00_000000000000", -- twrite, gr3
 385 => b"00000_0010_00_001010010101", -- load, gr2, P2BOMB4POS
 386 => b"00011_0010_01_000000000000", -- sub, gr2
 387 => b"00000_0000_00_000000001111", -- 15
 388 => b"10000_0010_00_000000000000", -- tpoint, gr2
 389 => b"01111_0000_00_000000000000", -- tread, gr0
 390 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 391 => b"00110_0000_01_000000000000", -- beq
 392 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 393 => b"01110_0011_00_000000000000", -- twrite, gr3
 394 => b"00011_0010_01_000000000000", -- sub, gr2
 395 => b"00000_0000_00_000000001111", -- 15
 396 => b"10000_0010_00_000000000000", -- tpoint, gr2
 397 => b"01111_0000_00_000000000000", -- tread, gr0
 398 => b"00011_0000_00_001010110010", -- sub, gr0, WALL
 399 => b"00110_0000_01_000000000000", -- beq
 400 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 401 => b"01110_0011_00_000000000000", -- twrite, gr3
 402 => b"00100_0000_01_000000000000", -- jump
 403 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 404 => b"10101_0000_01_000000000000", -- btn1
 405 => b"00000_0000_00_000110011010", -- BTN1
 406 => b"11010_0000_01_000000000000", -- btn2
 407 => b"00000_0000_00_000110111111", -- BTN2
 408 => b"00100_0000_01_000000000000", -- jump
 409 => b"00000_0000_00_000000000100", -- BUTTON_R
 410 => b"00000_0000_00_001010100111", -- load, gr0, P1BOMBCOUNT
 411 => b"00011_0000_00_001010101001", -- sub, gr0, MAXBOMBS
 412 => b"00110_0000_01_000000000000", -- beq
 413 => b"00000_0000_00_000110010110", -- BTN1_R
 414 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 415 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 416 => b"00000_0000_00_001010101011", -- load, gr0, YPOS1
 417 => b"01000_0000_01_000000000000", -- mul, gr0
 418 => b"00000_0000_00_000000001111", -- 15
 419 => b"00010_0000_00_001010101010", -- add, gr0, XPOS1
 420 => b"10000_0000_00_000000000000", -- tpoint, gr0
 421 => b"01111_0001_00_000000000000", -- tread, gr1
 422 => b"00011_0001_00_001010110101", -- sub, gr1, EGG
 423 => b"00110_0000_01_000000000000", -- beq
 424 => b"00000_0000_00_000110010110", -- BTN1_R
 425 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 426 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 427 => b"00000_0011_00_001010101011", -- load, gr3, YPOS1
 428 => b"00000_0010_00_001010110101", -- load, gr2, EGG
 429 => b"01000_0011_01_000000000000", -- mul, gr3
 430 => b"00000_0000_00_000000001111", -- 15
 431 => b"00010_0011_00_001010101010", -- add, gr3, XPOS1
 432 => b"10000_0011_00_000000000000", -- tpoint, gr3
 433 => b"01110_0010_00_000000000000", -- twrite, gr2
 434 => b"00000_0000_01_000000000000", -- load, gr0
 435 => b"00000_0000_00_000000000001", -- 1
 436 => b"00001_0000_10_001010000101", -- store, gr0, P1BOMB1ACTIVE
 437 => b"00001_0011_10_001010000011", -- store, gr3, P1BOMB1POS
 438 => b"00000_0000_01_000000000000", -- load, gr0
 439 => b"00000_0000_00_000000010000", -- 16
 440 => b"00001_0000_10_001010000100", -- store, gr0, P1BOMB1TIME
 441 => b"00000_0000_00_001010100111", -- load, gr0, P1BOMBCOUNT
 442 => b"00010_0000_01_000000000000", -- add, gr0
 443 => b"00000_0000_00_000000000001", -- 1
 444 => b"00001_0000_10_001010100111", -- store, gr0, P1BOMBCOUNT
 445 => b"00100_0000_01_000000000000", -- jump
 446 => b"00000_0000_00_000110010110", -- BTN1_R
 447 => b"00000_0000_00_001010101000", -- load, gr0, P2BOMBCOUNT
 448 => b"00011_0000_00_001010101001", -- sub, gr0, MAXBOMBS
 449 => b"00110_0000_01_000000000000", -- beq
 450 => b"00000_0000_00_000110011000", -- BTN2_R
 451 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 452 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 453 => b"00000_0000_00_001010101101", -- load, gr0, YPOS2
 454 => b"01000_0000_01_000000000000", -- mul, gr0
 455 => b"00000_0000_00_000000001111", -- 15
 456 => b"00010_0000_00_001010101100", -- add, gr0, XPOS2
 457 => b"10000_0000_00_000000000000", -- tpoint, gr0
 458 => b"01111_0001_00_000000000000", -- tread, gr1
 459 => b"00011_0001_00_001010110101", -- sub, gr1, EGG
 460 => b"00110_0000_01_000000000000", -- beq
 461 => b"00000_0000_00_000110011000", -- BTN2_R
 462 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 463 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 464 => b"00000_0011_00_001010101101", -- load, gr3, YPOS2
 465 => b"00000_0010_00_001010110101", -- load, gr2, EGG
 466 => b"01000_0011_01_000000000000", -- mul, gr3
 467 => b"00000_0000_00_000000001111", -- 15
 468 => b"00010_0011_00_001010101100", -- add, gr3, XPOS2
 469 => b"10000_0011_00_000000000000", -- tpoint, gr3
 470 => b"01110_0010_00_000000000000", -- twrite, gr2
 471 => b"00000_0000_01_000000000000", -- load, gr0
 472 => b"00000_0000_00_000000000001", -- 1
 473 => b"00001_0000_10_001010010111", -- store, gr0, P2BOMB4ACTIVE
 474 => b"00001_0011_10_001010010101", -- store, gr3, P2BOMB4POS
 475 => b"00000_0000_01_000000000000", -- load, gr0
 476 => b"00000_0000_00_000000010000", -- 16
 477 => b"00001_0000_10_001010010110", -- store, gr0, P2BOMB4TIME
 478 => b"00000_0000_00_001010101000", -- load, gr0, P2BOMBCOUNT
 479 => b"00010_0000_01_000000000000", -- add, gr0
 480 => b"00000_0000_00_000000000001", -- 1
 481 => b"00001_0000_10_001010101000", -- store, gr0, P2BOMBCOUNT
 482 => b"00100_0000_01_000000000000", -- jump
 483 => b"00000_0000_00_000110011000", -- BTN2_R
 484 => b"00000_0000_00_000000000000", -- 0
 485 => b"00100_0000_01_000000000000", -- jump
 486 => b"00000_0000_00_001010000001", -- COUNT1
 487 => b"10001_0000_01_000000000000", -- joy1r
 488 => b"00000_0000_00_000111111001", -- P1R
 489 => b"10011_0000_01_000000000000", -- joy1l
 490 => b"00000_0000_00_001000011011", -- P1L
 491 => b"10010_0000_01_000000000000", -- joy1u
 492 => b"00000_0000_00_001000001010", -- P1U
 493 => b"10100_0000_01_000000000000", -- joy1d
 494 => b"00000_0000_00_001000101100", -- P1D
 495 => b"10110_0000_01_000000000000", -- joy2r
 496 => b"00000_0000_00_001000111101", -- P2R
 497 => b"11000_0000_01_000000000000", -- joy2l
 498 => b"00000_0000_00_001001011111", -- P2L
 499 => b"10111_0000_01_000000000000", -- joy2u
 500 => b"00000_0000_00_001001001110", -- P2U
 501 => b"11001_0000_01_000000000000", -- joy2d
 502 => b"00000_0000_00_001001110000", -- P2D
 503 => b"00100_0000_01_000000000000", -- jump
 504 => b"00000_0000_00_000000000010", -- CONTROL_R
 505 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 506 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 507 => b"00000_0000_00_001010101011", -- load, gr0, YPOS1
 508 => b"01000_0000_01_000000000000", -- mul, gr0
 509 => b"00000_0000_00_000000001111", -- 15
 510 => b"00010_0000_00_001010101010", -- add, gr0, XPOS1
 511 => b"00010_0000_01_000000000000", -- add, gr0
 512 => b"00000_0000_00_000000000001", -- 1
 513 => b"10000_0000_00_000000000000", -- tpoint, gr0
 514 => b"01111_0001_00_000000000000", -- tread, gr1
 515 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 516 => b"00111_0000_01_000000000000", -- bne
 517 => b"00000_0000_00_000111101011", -- J1
 518 => b"00010_1100_01_000000000000", -- add, gr12
 519 => b"00000_0000_00_000000000001", -- 1
 520 => b"00100_0000_01_000000000000", -- jump
 521 => b"00000_0000_00_000111101011", -- J1
 522 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 523 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 524 => b"00000_0000_00_001010101011", -- load, gr0, YPOS1
 525 => b"00011_0000_01_000000000000", -- sub, gr0
 526 => b"00000_0000_00_000000000001", -- 1
 527 => b"01000_0000_01_000000000000", -- mul, gr0
 528 => b"00000_0000_00_000000001111", -- 15
 529 => b"00010_0000_00_001010101010", -- add, gr0, XPOS1
 530 => b"10000_0000_00_000000000000", -- tpoint, gr0
 531 => b"01111_0001_00_000000000000", -- tread, gr1
 532 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 533 => b"00111_0000_01_000000000000", -- bne
 534 => b"00000_0000_00_000111101111", -- J2
 535 => b"00011_1101_01_000000000000", -- sub, gr13
 536 => b"00000_0000_00_000000000001", -- 1
 537 => b"00100_0000_01_000000000000", -- jump
 538 => b"00000_0000_00_000111101111", -- J2
 539 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 540 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 541 => b"00000_0000_00_001010101011", -- load, gr0, YPOS1
 542 => b"01000_0000_01_000000000000", -- mul, gr0
 543 => b"00000_0000_00_000000001111", -- 15
 544 => b"00010_0000_00_001010101010", -- add, gr0, XPOS1
 545 => b"00011_0000_01_000000000000", -- sub, gr0
 546 => b"00000_0000_00_000000000001", -- 1
 547 => b"10000_0000_00_000000000000", -- tpoint, gr0
 548 => b"01111_0001_00_000000000000", -- tread, gr1
 549 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 550 => b"00111_0000_01_000000000000", -- bne
 551 => b"00000_0000_00_000111101011", -- J1
 552 => b"00011_1100_01_000000000000", -- sub, gr12
 553 => b"00000_0000_00_000000000001", -- 1
 554 => b"00100_0000_01_000000000000", -- jump
 555 => b"00000_0000_00_000111101011", -- J1
 556 => b"00001_1100_10_001010101010", -- store, gr12, XPOS1
 557 => b"00001_1101_10_001010101011", -- store, gr13, YPOS1
 558 => b"00000_0000_00_001010101011", -- load, gr0, YPOS1
 559 => b"00010_0000_01_000000000000", -- add, gr0
 560 => b"00000_0000_00_000000000001", -- 1
 561 => b"01000_0000_01_000000000000", -- mul, gr0
 562 => b"00000_0000_00_000000001111", -- 15
 563 => b"00010_0000_00_001010101010", -- add, gr0, XPOS1
 564 => b"10000_0000_00_000000000000", -- tpoint, gr0
 565 => b"01111_0001_00_000000000000", -- tread, gr1
 566 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 567 => b"00111_0000_01_000000000000", -- bne
 568 => b"00000_0000_00_000111101111", -- J2
 569 => b"00010_1101_01_000000000000", -- add, gr13
 570 => b"00000_0000_00_000000000001", -- 1
 571 => b"00100_0000_01_000000000000", -- jump
 572 => b"00000_0000_00_000111101111", -- J2
 573 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 574 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 575 => b"00000_0000_00_001010101101", -- load, gr0, YPOS2
 576 => b"01000_0000_01_000000000000", -- mul, gr0
 577 => b"00000_0000_00_000000001111", -- 15
 578 => b"00010_0000_00_001010101100", -- add, gr0, XPOS2
 579 => b"00010_0000_01_000000000000", -- add, gr0
 580 => b"00000_0000_00_000000000001", -- 1
 581 => b"10000_0000_00_000000000000", -- tpoint, gr0
 582 => b"01111_0001_00_000000000000", -- tread, gr1
 583 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 584 => b"00111_0000_01_000000000000", -- bne
 585 => b"00000_0000_00_000111110011", -- J3
 586 => b"00010_1110_01_000000000000", -- add, gr14
 587 => b"00000_0000_00_000000000001", -- 1
 588 => b"00100_0000_01_000000000000", -- jump
 589 => b"00000_0000_00_000111110011", -- J3
 590 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 591 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 592 => b"00000_0000_00_001010101101", -- load, gr0, YPOS2
 593 => b"00011_0000_01_000000000000", -- sub, gr0
 594 => b"00000_0000_00_000000000001", -- 1
 595 => b"01000_0000_01_000000000000", -- mul, gr0
 596 => b"00000_0000_00_000000001111", -- 15
 597 => b"00010_0000_00_001010101100", -- add, gr0, XPOS2
 598 => b"10000_0000_00_000000000000", -- tpoint, gr0
 599 => b"01111_0001_00_000000000000", -- tread, gr1
 600 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 601 => b"00111_0000_01_000000000000", -- bne
 602 => b"00000_0000_00_000000000010", -- CONTROL_R
 603 => b"00011_1111_01_000000000000", -- sub, gr15
 604 => b"00000_0000_00_000000000001", -- 1
 605 => b"00100_0000_01_000000000000", -- jump
 606 => b"00000_0000_00_000000000010", -- CONTROL_R
 607 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 608 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 609 => b"00000_0000_00_001010101101", -- load, gr0, YPOS2
 610 => b"01000_0000_01_000000000000", -- mul, gr0
 611 => b"00000_0000_00_000000001111", -- 15
 612 => b"00010_0000_00_001010101100", -- add, gr0, XPOS2
 613 => b"00011_0000_01_000000000000", -- sub, gr0
 614 => b"00000_0000_00_000000000001", -- 1
 615 => b"10000_0000_00_000000000000", -- tpoint, gr0
 616 => b"01111_0001_00_000000000000", -- tread, gr1
 617 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 618 => b"00111_0000_01_000000000000", -- bne
 619 => b"00000_0000_00_000111110011", -- J3
 620 => b"00011_1110_01_000000000000", -- sub, gr14
 621 => b"00000_0000_00_000000000001", -- 1
 622 => b"00100_0000_01_000000000000", -- jump
 623 => b"00000_0000_00_000111110011", -- J3
 624 => b"00001_1110_10_001010101100", -- store, gr14, XPOS2
 625 => b"00001_1111_10_001010101101", -- store, gr15, YPOS2
 626 => b"00000_0000_00_001010101101", -- load, gr0, YPOS2
 627 => b"00010_0000_01_000000000000", -- add, gr0
 628 => b"00000_0000_00_000000000001", -- 1
 629 => b"01000_0000_01_000000000000", -- mul, gr0
 630 => b"00000_0000_00_000000001111", -- 15
 631 => b"00010_0000_00_001010101100", -- add, gr0, XPOS2
 632 => b"10000_0000_00_000000000000", -- tpoint, gr0
 633 => b"01111_0001_00_000000000000", -- tread, gr1
 634 => b"00011_0001_00_001010110001", -- sub, gr1, GRASS
 635 => b"00111_0000_01_000000000000", -- bne
 636 => b"00000_0000_00_000000000010", -- CONTROL_R
 637 => b"00010_1111_01_000000000000", -- add, gr15
 638 => b"00000_0000_00_000000000001", -- 1
 639 => b"00100_0000_01_000000000000", -- jump
 640 => b"00000_0000_00_000000000010", -- CONTROL_R
 641 => b"00100_0000_01_000000000000", -- jump
 642 => b"00000_0000_00_000111100111", -- COUNT_R
 643 => b"00000_0000_00_000000000000", -- 0
 644 => b"00000_0000_00_000000000000", -- 0
 645 => b"00000_0000_00_000000000000", -- 0
 646 => b"00000_0000_00_000000000000", -- 0
 647 => b"00000_0000_00_000000000000", -- 0
 648 => b"00000_0000_00_000000000000", -- 0
 649 => b"00000_0000_00_000000000000", -- 0
 650 => b"00000_0000_00_000000000000", -- 0
 651 => b"00000_0000_00_000000000000", -- 0
 652 => b"00000_0000_00_000000000000", -- 0
 653 => b"00000_0000_00_000000000000", -- 0
 654 => b"00000_0000_00_000000000000", -- 0
 655 => b"00000_0000_00_000000000000", -- 0
 656 => b"00000_0000_00_000000000000", -- 0
 657 => b"00000_0000_00_000000000000", -- 0
 658 => b"00000_0000_00_000000000000", -- 0
 659 => b"00000_0000_00_000000000000", -- 0
 660 => b"00000_0000_00_000000000000", -- 0
 661 => b"00000_0000_00_000000000000", -- 0
 662 => b"00000_0000_00_000000000000", -- 0
 663 => b"00000_0000_00_000000000000", -- 0
 664 => b"00000_0000_00_000000000000", -- 0
 665 => b"00000_0000_00_000000000000", -- 0
 666 => b"00000_0000_00_000000000000", -- 0
 667 => b"00000_0000_00_000000000000", -- 0
 668 => b"00000_0000_00_000000000000", -- 0
 669 => b"00000_0000_00_000000000000", -- 0
 670 => b"00000_0000_00_000000000000", -- 0
 671 => b"00000_0000_00_000000000000", -- 0
 672 => b"00000_0000_00_000000000000", -- 0
 673 => b"00000_0000_00_000000000000", -- 0
 674 => b"00000_0000_00_000000000000", -- 0
 675 => b"00000_0000_00_000000000000", -- 0
 676 => b"00000_0000_00_000000000000", -- 0
 677 => b"00000_0000_00_000000000000", -- 0
 678 => b"00000_0000_00_000000000000", -- 0
 679 => b"00000_0000_00_000000000000", -- 0
 680 => b"00000_0000_00_000000000000", -- 0
 681 => b"00000_0000_00_000000000001", -- 1
 682 => b"00000_0000_00_000000000000", -- 0
 683 => b"00000_0000_00_000000000000", -- 0
 684 => b"00000_0000_00_000000000000", -- 0
 685 => b"00000_0000_00_000000000000", -- 0
 686 => b"00000_0000_00_000000000000", -- 0
 687 => b"00000_0000_00_000000000000", -- 0
 688 => b"00000_0000_00_000000000000", -- 0
 689 => b"00000_0000_00_000000000000", -- 0
 690 => b"00000_0000_00_000000000001", -- 1
 691 => b"00000_0000_00_000000000010", -- 2
 692 => b"00000_0000_00_000000000011", -- 3
 693 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
