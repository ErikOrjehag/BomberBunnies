library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_001001111101", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000111000011", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011000100", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000010000", -- BOOM1
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000001101010", -- BOOM2
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  16 => b"00000_0000_00_001100011111", -- load, gr0, P1EXPLOSION1ACTIVE
  17 => b"00011_0000_01_000000000000", -- sub, gr0
  18 => b"00000_0000_00_000000000001", -- 1
  19 => b"00111_0000_01_000000000000", -- bne
  20 => b"00000_0000_00_000000001100", -- BOOM1_R
  21 => b"00000_0000_00_001100011110", -- load, gr0, P1EXPLOSION1TIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000001", -- 1
  24 => b"00001_0000_10_001100011110", -- store, gr0, P1EXPLOSION1TIME
  25 => b"00000_0000_00_001100011110", -- load, gr0, P1EXPLOSION1TIME
  26 => b"00011_0000_01_000000000000", -- sub, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00111_0000_01_000000000000", -- bne
  29 => b"00000_0000_00_000000001100", -- BOOM1_R
  30 => b"00000_0000_01_000000000000", -- load, gr0
  31 => b"00000_0000_00_000000000000", -- 0
  32 => b"00001_0000_10_001100011111", -- store, gr0, P1EXPLOSION1ACTIVE
  33 => b"00000_0010_00_001100100000", -- load, gr2, P1EXPLOSION1POS
  34 => b"00000_0011_00_001101001001", -- load, gr3, GRASS
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01110_0011_00_000000000000", -- twrite, gr3
  37 => b"00010_0010_01_000000000000", -- add, gr2
  38 => b"00000_0000_00_000000000001", -- 1
  39 => b"10000_0010_00_000000000000", -- tpoint, gr2
  40 => b"01111_0000_00_000000000000", -- tread, gr0
  41 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  42 => b"00111_0000_01_000000000000", -- bne
  43 => b"00000_0000_00_000000110101", -- E1LEFT
  44 => b"01110_0011_00_000000000000", -- twrite, gr3
  45 => b"00010_0010_01_000000000000", -- add, gr2
  46 => b"00000_0000_00_000000000001", -- 1
  47 => b"10000_0010_00_000000000000", -- tpoint, gr2
  48 => b"01111_0000_00_000000000000", -- tread, gr0
  49 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  50 => b"00111_0000_01_000000000000", -- bne
  51 => b"00000_0000_00_000000110101", -- E1LEFT
  52 => b"01110_0011_00_000000000000", -- twrite, gr3
  53 => b"00000_0010_00_001100100000", -- load, gr2, P1EXPLOSION1POS
  54 => b"00011_0010_01_000000000000", -- sub, gr2
  55 => b"00000_0000_00_000000000001", -- 1
  56 => b"10000_0010_00_000000000000", -- tpoint, gr2
  57 => b"01111_0000_00_000000000000", -- tread, gr0
  58 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  59 => b"00111_0000_01_000000000000", -- bne
  60 => b"00000_0000_00_000001000110", -- E1DOWN
  61 => b"01110_0011_00_000000000000", -- twrite, gr3
  62 => b"00011_0010_01_000000000000", -- sub, gr2
  63 => b"00000_0000_00_000000000001", -- 1
  64 => b"10000_0010_00_000000000000", -- tpoint, gr2
  65 => b"01111_0000_00_000000000000", -- tread, gr0
  66 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  67 => b"00111_0000_01_000000000000", -- bne
  68 => b"00000_0000_00_000001000110", -- E1DOWN
  69 => b"01110_0011_00_000000000000", -- twrite, gr3
  70 => b"00000_0010_00_001100100000", -- load, gr2, P1EXPLOSION1POS
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000001111", -- 15
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0000_00_000000000000", -- tread, gr0
  75 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  76 => b"00111_0000_01_000000000000", -- bne
  77 => b"00000_0000_00_000001010111", -- E1UP
  78 => b"01110_0011_00_000000000000", -- twrite, gr3
  79 => b"00010_0010_01_000000000000", -- add, gr2
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"10000_0010_00_000000000000", -- tpoint, gr2
  82 => b"01111_0000_00_000000000000", -- tread, gr0
  83 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  84 => b"00111_0000_01_000000000000", -- bne
  85 => b"00000_0000_00_000001010111", -- E1UP
  86 => b"01110_0011_00_000000000000", -- twrite, gr3
  87 => b"00000_0010_00_001100100000", -- load, gr2, P1EXPLOSION1POS
  88 => b"00011_0010_01_000000000000", -- sub, gr2
  89 => b"00000_0000_00_000000001111", -- 15
  90 => b"10000_0010_00_000000000000", -- tpoint, gr2
  91 => b"01111_0000_00_000000000000", -- tread, gr0
  92 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
  93 => b"00111_0000_01_000000000000", -- bne
  94 => b"00000_0000_00_000000001100", -- BOOM1_R
  95 => b"01110_0011_00_000000000000", -- twrite, gr3
  96 => b"00011_0010_01_000000000000", -- sub, gr2
  97 => b"00000_0000_00_000000001111", -- 15
  98 => b"10000_0010_00_000000000000", -- tpoint, gr2
  99 => b"01111_0000_00_000000000000", -- tread, gr0
 100 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 101 => b"00111_0000_01_000000000000", -- bne
 102 => b"00000_0000_00_000000001100", -- BOOM1_R
 103 => b"01110_0011_00_000000000000", -- twrite, gr3
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000000001100", -- BOOM1_R
 106 => b"00000_0000_00_001100110001", -- load, gr0, P2EXPLOSION1ACTIVE
 107 => b"00011_0000_01_000000000000", -- sub, gr0
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00111_0000_01_000000000000", -- bne
 110 => b"00000_0000_00_000000001110", -- BOOM2_R
 111 => b"00000_0000_00_001100110000", -- load, gr0, P2EXPLOSION1TIME
 112 => b"00011_0000_01_000000000000", -- sub, gr0
 113 => b"00000_0000_00_000000000001", -- 1
 114 => b"00001_0000_10_001100110000", -- store, gr0, P2EXPLOSION1TIME
 115 => b"00000_0000_00_001100110000", -- load, gr0, P2EXPLOSION1TIME
 116 => b"00011_0000_01_000000000000", -- sub, gr0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00111_0000_01_000000000000", -- bne
 119 => b"00000_0000_00_000000001110", -- BOOM2_R
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001100110001", -- store, gr0, P2EXPLOSION1ACTIVE
 123 => b"00000_0010_00_001100110010", -- load, gr2, P2EXPLOSION1POS
 124 => b"00000_0011_00_001101001001", -- load, gr3, GRASS
 125 => b"10000_0010_00_000000000000", -- tpoint, gr2
 126 => b"01110_0011_00_000000000000", -- twrite, gr3
 127 => b"00010_0010_01_000000000000", -- add, gr2
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"10000_0010_00_000000000000", -- tpoint, gr2
 130 => b"01111_0000_00_000000000000", -- tread, gr0
 131 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 132 => b"00111_0000_01_000000000000", -- bne
 133 => b"00000_0000_00_000010001111", -- E2LEFT
 134 => b"01110_0011_00_000000000000", -- twrite, gr3
 135 => b"00010_0010_01_000000000000", -- add, gr2
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0010_00_000000000000", -- tpoint, gr2
 138 => b"01111_0000_00_000000000000", -- tread, gr0
 139 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000010001111", -- E2LEFT
 142 => b"01110_0011_00_000000000000", -- twrite, gr3
 143 => b"00000_0010_00_001100110010", -- load, gr2, P2EXPLOSION1POS
 144 => b"00011_0010_01_000000000000", -- sub, gr2
 145 => b"00000_0000_00_000000000001", -- 1
 146 => b"10000_0010_00_000000000000", -- tpoint, gr2
 147 => b"01111_0000_00_000000000000", -- tread, gr0
 148 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 149 => b"00111_0000_01_000000000000", -- bne
 150 => b"00000_0000_00_000010100000", -- E2DOWN
 151 => b"01110_0011_00_000000000000", -- twrite, gr3
 152 => b"00011_0010_01_000000000000", -- sub, gr2
 153 => b"00000_0000_00_000000000001", -- 1
 154 => b"10000_0010_00_000000000000", -- tpoint, gr2
 155 => b"01111_0000_00_000000000000", -- tread, gr0
 156 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000010100000", -- E2DOWN
 159 => b"01110_0011_00_000000000000", -- twrite, gr3
 160 => b"00000_0010_00_001100110010", -- load, gr2, P2EXPLOSION1POS
 161 => b"00010_0010_01_000000000000", -- add, gr2
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"10000_0010_00_000000000000", -- tpoint, gr2
 164 => b"01111_0000_00_000000000000", -- tread, gr0
 165 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 166 => b"00111_0000_01_000000000000", -- bne
 167 => b"00000_0000_00_000010110001", -- E2UP
 168 => b"01110_0011_00_000000000000", -- twrite, gr3
 169 => b"00010_0010_01_000000000000", -- add, gr2
 170 => b"00000_0000_00_000000001111", -- 15
 171 => b"10000_0010_00_000000000000", -- tpoint, gr2
 172 => b"01111_0000_00_000000000000", -- tread, gr0
 173 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000010110001", -- E2UP
 176 => b"01110_0011_00_000000000000", -- twrite, gr3
 177 => b"00000_0010_00_001100110010", -- load, gr2, P2EXPLOSION1POS
 178 => b"00011_0010_01_000000000000", -- sub, gr2
 179 => b"00000_0000_00_000000001111", -- 15
 180 => b"10000_0010_00_000000000000", -- tpoint, gr2
 181 => b"01111_0000_00_000000000000", -- tread, gr0
 182 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 183 => b"00111_0000_01_000000000000", -- bne
 184 => b"00000_0000_00_000000001110", -- BOOM2_R
 185 => b"01110_0011_00_000000000000", -- twrite, gr3
 186 => b"00011_0010_01_000000000000", -- sub, gr2
 187 => b"00000_0000_00_000000001111", -- 15
 188 => b"10000_0010_00_000000000000", -- tpoint, gr2
 189 => b"01111_0000_00_000000000000", -- tread, gr0
 190 => b"00011_0000_00_001101001100", -- sub, gr0, EXPLOSION
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000001110", -- BOOM2_R
 193 => b"01110_0011_00_000000000000", -- twrite, gr3
 194 => b"00100_0000_01_000000000000", -- jump
 195 => b"00000_0000_00_000000001110", -- BOOM2_R
 196 => b"00000_0000_00_001100011101", -- load, gr0, P1BOMB1ACTIVE
 197 => b"00011_0000_01_000000000000", -- sub, gr0
 198 => b"00000_0000_00_000000000001", -- 1
 199 => b"00111_0000_01_000000000000", -- bne
 200 => b"00000_0000_00_000011010010", -- P1BOMB2
 201 => b"00000_0000_00_001100011100", -- load, gr0, P1BOMB1TIME
 202 => b"00011_0000_01_000000000000", -- sub, gr0
 203 => b"00000_0000_00_000000000001", -- 1
 204 => b"00001_0000_10_001100011100", -- store, gr0, P1BOMB1TIME
 205 => b"00000_0000_01_000000000000", -- load, gr0
 206 => b"00000_0000_00_000000000000", -- 0
 207 => b"00011_0000_00_001100011100", -- sub, gr0, P1BOMB1TIME
 208 => b"00110_0000_01_000000000000", -- beq
 209 => b"00000_0000_00_000100011100", -- P1EXPLOSION1INIT
 210 => b"00000_0000_00_001100100011", -- load, gr0, P1BOMB2ACTIVE
 211 => b"00011_0000_01_000000000000", -- sub, gr0
 212 => b"00000_0000_00_000000000001", -- 1
 213 => b"00111_0000_01_000000000000", -- bne
 214 => b"00000_0000_00_000011100000", -- P1BOMB3
 215 => b"00000_0000_00_001100100010", -- load, gr0, P1BOMB2TIME
 216 => b"00011_0000_01_000000000000", -- sub, gr0
 217 => b"00000_0000_00_000000000001", -- 1
 218 => b"00001_0000_10_001100100010", -- store, gr0, P1BOMB2TIME
 219 => b"00000_0000_01_000000000000", -- load, gr0
 220 => b"00000_0000_00_000000000000", -- 0
 221 => b"00011_0000_00_001100100010", -- sub, gr0, P1BOMB2TIME
 222 => b"00110_0000_01_000000000000", -- beq
 223 => b"00000_0000_00_000100101011", -- P1EXPLOSION2INIT
 224 => b"00000_0000_00_001100101001", -- load, gr0, P1BOMB3ACTIVE
 225 => b"00011_0000_01_000000000000", -- sub, gr0
 226 => b"00000_0000_00_000000000001", -- 1
 227 => b"00111_0000_01_000000000000", -- bne
 228 => b"00000_0000_00_000011110000", -- P2BOMB1
 229 => b"00000_0000_00_001100101000", -- load, gr0, P1BOMB3TIME
 230 => b"00011_0000_01_000000000000", -- sub, gr0
 231 => b"00000_0000_00_000000000001", -- 1
 232 => b"00001_0000_10_001100101000", -- store, gr0, P1BOMB3TIME
 233 => b"00000_0000_01_000000000000", -- load, gr0
 234 => b"00000_0000_00_000000000000", -- 0
 235 => b"00011_0000_00_001100101000", -- sub, gr0, P1BOMB3TIME
 236 => b"00110_0000_01_000000000000", -- beq
 237 => b"00000_0000_00_000100111010", -- P1EXPLOSION3INIT
 238 => b"00100_0000_01_000000000000", -- jump
 239 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 240 => b"00000_0000_00_001100101111", -- load, gr0, P2BOMB1ACTIVE
 241 => b"00011_0000_01_000000000000", -- sub, gr0
 242 => b"00000_0000_00_000000000001", -- 1
 243 => b"00111_0000_01_000000000000", -- bne
 244 => b"00000_0000_00_000011111110", -- P2BOMB2
 245 => b"00000_0000_00_001100101110", -- load, gr0, P2BOMB1TIME
 246 => b"00011_0000_01_000000000000", -- sub, gr0
 247 => b"00000_0000_00_000000000001", -- 1
 248 => b"00001_0000_10_001100101110", -- store, gr0, P2BOMB1TIME
 249 => b"00000_0000_01_000000000000", -- load, gr0
 250 => b"00000_0000_00_000000000000", -- 0
 251 => b"00011_0000_00_001100101110", -- sub, gr0, P2BOMB1TIME
 252 => b"00110_0000_01_000000000000", -- beq
 253 => b"00000_0000_00_000101001001", -- P2EXPLOSION1INIT
 254 => b"00000_0000_00_001100110101", -- load, gr0, P2BOMB2ACTIVE
 255 => b"00011_0000_01_000000000000", -- sub, gr0
 256 => b"00000_0000_00_000000000001", -- 1
 257 => b"00111_0000_01_000000000000", -- bne
 258 => b"00000_0000_00_000100001100", -- P2BOMB3
 259 => b"00000_0000_00_001100110100", -- load, gr0, P2BOMB2TIME
 260 => b"00011_0000_01_000000000000", -- sub, gr0
 261 => b"00000_0000_00_000000000001", -- 1
 262 => b"00001_0000_10_001100110100", -- store, gr0, P2BOMB2TIME
 263 => b"00000_0000_01_000000000000", -- load, gr0
 264 => b"00000_0000_00_000000000000", -- 0
 265 => b"00011_0000_00_001100110100", -- sub, gr0, P2BOMB2TIME
 266 => b"00110_0000_01_000000000000", -- beq
 267 => b"00000_0000_00_000101011000", -- P2EXPLOSION2INIT
 268 => b"00000_0000_00_001100111011", -- load, gr0, P2BOMB3ACTIVE
 269 => b"00011_0000_01_000000000000", -- sub, gr0
 270 => b"00000_0000_00_000000000001", -- 1
 271 => b"00111_0000_01_000000000000", -- bne
 272 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 273 => b"00000_0000_00_001100111010", -- load, gr0, P2BOMB3TIME
 274 => b"00011_0000_01_000000000000", -- sub, gr0
 275 => b"00000_0000_00_000000000001", -- 1
 276 => b"00001_0000_10_001100111010", -- store, gr0, P2BOMB3TIME
 277 => b"00000_0000_01_000000000000", -- load, gr0
 278 => b"00000_0000_00_000000000000", -- 0
 279 => b"00011_0000_00_001100111010", -- sub, gr0, P2BOMB3TIME
 280 => b"00110_0000_01_000000000000", -- beq
 281 => b"00000_0000_00_000101100111", -- P2EXPLOSION3INIT
 282 => b"00100_0000_01_000000000000", -- jump
 283 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 284 => b"00000_0000_00_001100011011", -- load, gr0, P1BOMB1POS
 285 => b"00001_0000_10_001100100000", -- store, gr0, P1EXPLOSION1POS
 286 => b"00000_0000_01_000000000000", -- load, gr0
 287 => b"00000_0000_00_000000000001", -- 1
 288 => b"00001_0000_10_001100011111", -- store, gr0, P1EXPLOSION1ACTIVE
 289 => b"00000_0000_01_000000000000", -- load, gr0
 290 => b"00000_0000_00_000000000010", -- 2
 291 => b"00001_0000_10_001100011110", -- store, gr0, P1EXPLOSION1TIME
 292 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 293 => b"00011_0000_01_000000000000", -- sub, gr0
 294 => b"00000_0000_00_000000000001", -- 1
 295 => b"00001_0000_10_001100111111", -- store, gr0, P1BOMBCOUNT
 296 => b"00000_0100_00_001100011011", -- load, gr4, P1BOMB1POS
 297 => b"00100_0000_01_000000000000", -- jump
 298 => b"00000_0000_00_000101110110", -- EXPLODE
 299 => b"00000_0000_00_001100100001", -- load, gr0, P1BOMB2POS
 300 => b"00001_0000_10_001100100110", -- store, gr0, P1EXPLOSION2POS
 301 => b"00000_0000_01_000000000000", -- load, gr0
 302 => b"00000_0000_00_000000000001", -- 1
 303 => b"00001_0000_10_001100100101", -- store, gr0, P1EXPLOSION2ACTIVE
 304 => b"00000_0000_01_000000000000", -- load, gr0
 305 => b"00000_0000_00_000000000010", -- 2
 306 => b"00001_0000_10_001100100100", -- store, gr0, P1EXPLOSION2TIME
 307 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 308 => b"00011_0000_01_000000000000", -- sub, gr0
 309 => b"00000_0000_00_000000000001", -- 1
 310 => b"00001_0000_10_001100111111", -- store, gr0, P1BOMBCOUNT
 311 => b"00000_0100_00_001100100001", -- load, gr4, P1BOMB2POS
 312 => b"00100_0000_01_000000000000", -- jump
 313 => b"00000_0000_00_000101110110", -- EXPLODE
 314 => b"00000_0000_00_001100100111", -- load, gr0, P1BOMB3POS
 315 => b"00001_0000_10_001100101100", -- store, gr0, P1EXPLOSION3POS
 316 => b"00000_0000_01_000000000000", -- load, gr0
 317 => b"00000_0000_00_000000000001", -- 1
 318 => b"00001_0000_10_001100101011", -- store, gr0, P1EXPLOSION3ACTIVE
 319 => b"00000_0000_01_000000000000", -- load, gr0
 320 => b"00000_0000_00_000000000010", -- 2
 321 => b"00001_0000_10_001100101010", -- store, gr0, P1EXPLOSION3TIME
 322 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 323 => b"00011_0000_01_000000000000", -- sub, gr0
 324 => b"00000_0000_00_000000000001", -- 1
 325 => b"00001_0000_10_001100111111", -- store, gr0, P1BOMBCOUNT
 326 => b"00000_0100_00_001100100111", -- load, gr4, P1BOMB3POS
 327 => b"00100_0000_01_000000000000", -- jump
 328 => b"00000_0000_00_000101110110", -- EXPLODE
 329 => b"00000_0000_00_001100101101", -- load, gr0, P2BOMB1POS
 330 => b"00001_0000_10_001100110010", -- store, gr0, P2EXPLOSION1POS
 331 => b"00000_0000_01_000000000000", -- load, gr0
 332 => b"00000_0000_00_000000000001", -- 1
 333 => b"00001_0000_10_001100110001", -- store, gr0, P2EXPLOSION1ACTIVE
 334 => b"00000_0000_01_000000000000", -- load, gr0
 335 => b"00000_0000_00_000000000010", -- 2
 336 => b"00001_0000_10_001100110000", -- store, gr0, P2EXPLOSION1TIME
 337 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 338 => b"00011_0000_01_000000000000", -- sub, gr0
 339 => b"00000_0000_00_000000000001", -- 1
 340 => b"00001_0000_10_001101000000", -- store, gr0, P2BOMBCOUNT
 341 => b"00000_0100_00_001100101101", -- load, gr4, P2BOMB1POS
 342 => b"00100_0000_01_000000000000", -- jump
 343 => b"00000_0000_00_000101110110", -- EXPLODE
 344 => b"00000_0000_00_001100110011", -- load, gr0, P2BOMB2POS
 345 => b"00001_0000_10_001100111000", -- store, gr0, P2EXPLOSION2POS
 346 => b"00000_0000_01_000000000000", -- load, gr0
 347 => b"00000_0000_00_000000000001", -- 1
 348 => b"00001_0000_10_001100110111", -- store, gr0, P2EXPLOSION2ACTIVE
 349 => b"00000_0000_01_000000000000", -- load, gr0
 350 => b"00000_0000_00_000000000010", -- 2
 351 => b"00001_0000_10_001100110110", -- store, gr0, P2EXPLOSION2TIME
 352 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 353 => b"00011_0000_01_000000000000", -- sub, gr0
 354 => b"00000_0000_00_000000000001", -- 1
 355 => b"00001_0000_10_001101000000", -- store, gr0, P2BOMBCOUNT
 356 => b"00000_0100_00_001100110011", -- load, gr4, P2BOMB2POS
 357 => b"00100_0000_01_000000000000", -- jump
 358 => b"00000_0000_00_000101110110", -- EXPLODE
 359 => b"00000_0000_00_001100111001", -- load, gr0, P2BOMB3POS
 360 => b"00001_0000_10_001100111110", -- store, gr0, P2EXPLOSION3POS
 361 => b"00000_0000_01_000000000000", -- load, gr0
 362 => b"00000_0000_00_000000000001", -- 1
 363 => b"00001_0000_10_001100111101", -- store, gr0, P2EXPLOSION3ACTIVE
 364 => b"00000_0000_01_000000000000", -- load, gr0
 365 => b"00000_0000_00_000000000010", -- 2
 366 => b"00001_0000_10_001100111100", -- store, gr0, P2EXPLOSION3TIME
 367 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 368 => b"00011_0000_01_000000000000", -- sub, gr0
 369 => b"00000_0000_00_000000000001", -- 1
 370 => b"00001_0000_10_001101000000", -- store, gr0, P2BOMBCOUNT
 371 => b"00000_0100_00_001100111001", -- load, gr4, P2BOMB3POS
 372 => b"00100_0000_01_000000000000", -- jump
 373 => b"00000_0000_00_000101110110", -- EXPLODE
 374 => b"00001_0100_10_001101000110", -- store, gr4, MOVE
 375 => b"00000_0010_00_001101000110", -- load, gr2, MOVE
 376 => b"00000_0011_00_001101001100", -- load, gr3, EXPLOSION
 377 => b"10000_0010_00_000000000000", -- tpoint, gr2
 378 => b"01110_0011_00_000000000000", -- twrite, gr3
 379 => b"00010_0010_01_000000000000", -- add, gr2
 380 => b"00000_0000_00_000000000001", -- 1
 381 => b"10000_0010_00_000000000000", -- tpoint, gr2
 382 => b"01111_0000_00_000000000000", -- tread, gr0
 383 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 384 => b"00110_0000_01_000000000000", -- beq
 385 => b"00000_0000_00_000110001011", -- EXPLODELEFT
 386 => b"01110_0011_00_000000000000", -- twrite, gr3
 387 => b"00010_0010_01_000000000000", -- add, gr2
 388 => b"00000_0000_00_000000000001", -- 1
 389 => b"10000_0010_00_000000000000", -- tpoint, gr2
 390 => b"01111_0000_00_000000000000", -- tread, gr0
 391 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 392 => b"00110_0000_01_000000000000", -- beq
 393 => b"00000_0000_00_000110001011", -- EXPLODELEFT
 394 => b"01110_0011_00_000000000000", -- twrite, gr3
 395 => b"00001_0100_10_001101000110", -- store, gr4, MOVE
 396 => b"00000_0010_00_001101000110", -- load, gr2, MOVE
 397 => b"00011_0010_01_000000000000", -- sub, gr2
 398 => b"00000_0000_00_000000000001", -- 1
 399 => b"10000_0010_00_000000000000", -- tpoint, gr2
 400 => b"01111_0000_00_000000000000", -- tread, gr0
 401 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 402 => b"00110_0000_01_000000000000", -- beq
 403 => b"00000_0000_00_000110011101", -- EXPLODEDOWN
 404 => b"01110_0011_00_000000000000", -- twrite, gr3
 405 => b"00011_0010_01_000000000000", -- sub, gr2
 406 => b"00000_0000_00_000000000001", -- 1
 407 => b"10000_0010_00_000000000000", -- tpoint, gr2
 408 => b"01111_0000_00_000000000000", -- tread, gr0
 409 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 410 => b"00110_0000_01_000000000000", -- beq
 411 => b"00000_0000_00_000110011101", -- EXPLODEDOWN
 412 => b"01110_0011_00_000000000000", -- twrite, gr3
 413 => b"00001_0100_10_001101000110", -- store, gr4, MOVE
 414 => b"00000_0010_00_001101000110", -- load, gr2, MOVE
 415 => b"00010_0010_01_000000000000", -- add, gr2
 416 => b"00000_0000_00_000000001111", -- 15
 417 => b"10000_0010_00_000000000000", -- tpoint, gr2
 418 => b"01111_0000_00_000000000000", -- tread, gr0
 419 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 420 => b"00110_0000_01_000000000000", -- beq
 421 => b"00000_0000_00_000110101111", -- EXPLODEUP
 422 => b"01110_0011_00_000000000000", -- twrite, gr3
 423 => b"00010_0010_01_000000000000", -- add, gr2
 424 => b"00000_0000_00_000000001111", -- 15
 425 => b"10000_0010_00_000000000000", -- tpoint, gr2
 426 => b"01111_0000_00_000000000000", -- tread, gr0
 427 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 428 => b"00110_0000_01_000000000000", -- beq
 429 => b"00000_0000_00_000110101111", -- EXPLODEUP
 430 => b"01110_0011_00_000000000000", -- twrite, gr3
 431 => b"00001_0100_10_001101000110", -- store, gr4, MOVE
 432 => b"00000_0010_00_001101000110", -- load, gr2, MOVE
 433 => b"00011_0010_01_000000000000", -- sub, gr2
 434 => b"00000_0000_00_000000001111", -- 15
 435 => b"10000_0010_00_000000000000", -- tpoint, gr2
 436 => b"01111_0000_00_000000000000", -- tread, gr0
 437 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 438 => b"00110_0000_01_000000000000", -- beq
 439 => b"00000_0000_00_000011000100", -- TICKBOMBS
 440 => b"01110_0011_00_000000000000", -- twrite, gr3
 441 => b"00011_0010_01_000000000000", -- sub, gr2
 442 => b"00000_0000_00_000000001111", -- 15
 443 => b"10000_0010_00_000000000000", -- tpoint, gr2
 444 => b"01111_0000_00_000000000000", -- tread, gr0
 445 => b"00011_0000_00_001101001010", -- sub, gr0, WALL
 446 => b"00110_0000_01_000000000000", -- beq
 447 => b"00000_0000_00_000011000100", -- TICKBOMBS
 448 => b"01110_0011_00_000000000000", -- twrite, gr3
 449 => b"00100_0000_01_000000000000", -- jump
 450 => b"00000_0000_00_000011000100", -- TICKBOMBS
 451 => b"10101_0000_01_000000000000", -- btn1
 452 => b"00000_0000_00_000111001001", -- BTN1
 453 => b"11010_0000_01_000000000000", -- btn2
 454 => b"00000_0000_00_001000100011", -- BTN2
 455 => b"00100_0000_01_000000000000", -- jump
 456 => b"00000_0000_00_000000000100", -- BUTTON_R
 457 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 458 => b"00011_0000_00_001101000001", -- sub, gr0, MAXBOMBS
 459 => b"00110_0000_01_000000000000", -- beq
 460 => b"00000_0000_00_000111000101", -- BTN1_R
 461 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 462 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 463 => b"00000_0000_00_001101000011", -- load, gr0, YPOS1
 464 => b"01000_0000_01_000000000000", -- mul, gr0
 465 => b"00000_0000_00_000000001111", -- 15
 466 => b"00010_0000_00_001101000010", -- add, gr0, XPOS1
 467 => b"10000_0000_00_000000000000", -- tpoint, gr0
 468 => b"01111_0001_00_000000000000", -- tread, gr1
 469 => b"00011_0001_00_001101001101", -- sub, gr1, EGG
 470 => b"00110_0000_01_000000000000", -- beq
 471 => b"00000_0000_00_000111000101", -- BTN1_R
 472 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 473 => b"00011_0000_01_000000000000", -- sub, gr0
 474 => b"00000_0000_00_000000000000", -- 0
 475 => b"00110_0000_01_000000000000", -- beq
 476 => b"00000_0000_00_000111101101", -- P1PLACEBOMB1
 477 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 478 => b"00011_0000_01_000000000000", -- sub, gr0
 479 => b"00000_0000_00_000000000001", -- 1
 480 => b"00110_0000_01_000000000000", -- beq
 481 => b"00000_0000_00_000111111111", -- P1PLACEBOMB2
 482 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 483 => b"00011_0000_01_000000000000", -- sub, gr0
 484 => b"00000_0000_00_000000000010", -- 2
 485 => b"00110_0000_01_000000000000", -- beq
 486 => b"00000_0000_00_001000010001", -- P1PLACEBOMB3
 487 => b"00000_0000_00_001100111111", -- load, gr0, P1BOMBCOUNT
 488 => b"00010_0000_01_000000000000", -- add, gr0
 489 => b"00000_0000_00_000000000001", -- 1
 490 => b"00001_0000_10_001100111111", -- store, gr0, P1BOMBCOUNT
 491 => b"00100_0000_01_000000000000", -- jump
 492 => b"00000_0000_00_000111000101", -- BTN1_R
 493 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 494 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 495 => b"00000_0011_00_001101000011", -- load, gr3, YPOS1
 496 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 497 => b"01000_0011_01_000000000000", -- mul, gr3
 498 => b"00000_0000_00_000000001111", -- 15
 499 => b"00010_0011_00_001101000010", -- add, gr3, XPOS1
 500 => b"10000_0011_00_000000000000", -- tpoint, gr3
 501 => b"01110_0010_00_000000000000", -- twrite, gr2
 502 => b"00000_0000_01_000000000000", -- load, gr0
 503 => b"00000_0000_00_000000000001", -- 1
 504 => b"00001_0000_10_001100011101", -- store, gr0, P1BOMB1ACTIVE
 505 => b"00001_0011_10_001100011011", -- store, gr3, P1BOMB1POS
 506 => b"00000_0000_01_000000000000", -- load, gr0
 507 => b"00000_0000_00_000000010000", -- 16
 508 => b"00001_0000_10_001100011100", -- store, gr0, P1BOMB1TIME
 509 => b"00100_0000_01_000000000000", -- jump
 510 => b"00000_0000_00_000111100111", -- P1INCREASEBOMBCOUNTER
 511 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 512 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 513 => b"00000_0011_00_001101000011", -- load, gr3, YPOS1
 514 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 515 => b"01000_0011_01_000000000000", -- mul, gr3
 516 => b"00000_0000_00_000000001111", -- 15
 517 => b"00010_0011_00_001101000010", -- add, gr3, XPOS1
 518 => b"10000_0011_00_000000000000", -- tpoint, gr3
 519 => b"01110_0010_00_000000000000", -- twrite, gr2
 520 => b"00000_0000_01_000000000000", -- load, gr0
 521 => b"00000_0000_00_000000000001", -- 1
 522 => b"00001_0000_10_001100100011", -- store, gr0, P1BOMB2ACTIVE
 523 => b"00001_0011_10_001100100001", -- store, gr3, P1BOMB2POS
 524 => b"00000_0000_01_000000000000", -- load, gr0
 525 => b"00000_0000_00_000000010000", -- 16
 526 => b"00001_0000_10_001100100010", -- store, gr0, P1BOMB2TIME
 527 => b"00100_0000_01_000000000000", -- jump
 528 => b"00000_0000_00_000111100111", -- P1INCREASEBOMBCOUNTER
 529 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 530 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 531 => b"00000_0011_00_001101000011", -- load, gr3, YPOS1
 532 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 533 => b"01000_0011_01_000000000000", -- mul, gr3
 534 => b"00000_0000_00_000000001111", -- 15
 535 => b"00010_0011_00_001101000010", -- add, gr3, XPOS1
 536 => b"10000_0011_00_000000000000", -- tpoint, gr3
 537 => b"01110_0010_00_000000000000", -- twrite, gr2
 538 => b"00000_0000_01_000000000000", -- load, gr0
 539 => b"00000_0000_00_000000000001", -- 1
 540 => b"00001_0000_10_001100101001", -- store, gr0, P1BOMB3ACTIVE
 541 => b"00001_0011_10_001100100111", -- store, gr3, P1BOMB3POS
 542 => b"00000_0000_01_000000000000", -- load, gr0
 543 => b"00000_0000_00_000000010000", -- 16
 544 => b"00001_0000_10_001100101000", -- store, gr0, P1BOMB3TIME
 545 => b"00100_0000_01_000000000000", -- jump
 546 => b"00000_0000_00_000111100111", -- P1INCREASEBOMBCOUNTER
 547 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 548 => b"00011_0000_00_001101000001", -- sub, gr0, MAXBOMBS
 549 => b"00110_0000_01_000000000000", -- beq
 550 => b"00000_0000_00_000111000111", -- BTN2_R
 551 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 552 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 553 => b"00000_0000_00_001101000101", -- load, gr0, YPOS2
 554 => b"01000_0000_01_000000000000", -- mul, gr0
 555 => b"00000_0000_00_000000001111", -- 15
 556 => b"00010_0000_00_001101000100", -- add, gr0, XPOS2
 557 => b"10000_0000_00_000000000000", -- tpoint, gr0
 558 => b"01111_0001_00_000000000000", -- tread, gr1
 559 => b"00011_0001_00_001101001101", -- sub, gr1, EGG
 560 => b"00110_0000_01_000000000000", -- beq
 561 => b"00000_0000_00_000111000111", -- BTN2_R
 562 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 563 => b"00011_0000_01_000000000000", -- sub, gr0
 564 => b"00000_0000_00_000000000000", -- 0
 565 => b"00110_0000_01_000000000000", -- beq
 566 => b"00000_0000_00_001001000111", -- P2PLACEBOMB1
 567 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 568 => b"00011_0000_01_000000000000", -- sub, gr0
 569 => b"00000_0000_00_000000000001", -- 1
 570 => b"00110_0000_01_000000000000", -- beq
 571 => b"00000_0000_00_001001011001", -- P2PLACEBOMB2
 572 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 573 => b"00011_0000_01_000000000000", -- sub, gr0
 574 => b"00000_0000_00_000000000010", -- 2
 575 => b"00110_0000_01_000000000000", -- beq
 576 => b"00000_0000_00_001001101011", -- P2PLACEBOMB3
 577 => b"00000_0000_00_001101000000", -- load, gr0, P2BOMBCOUNT
 578 => b"00010_0000_01_000000000000", -- add, gr0
 579 => b"00000_0000_00_000000000001", -- 1
 580 => b"00001_0000_10_001101000000", -- store, gr0, P2BOMBCOUNT
 581 => b"00100_0000_01_000000000000", -- jump
 582 => b"00000_0000_00_000111000111", -- BTN2_R
 583 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 584 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 585 => b"00000_0011_00_001101000101", -- load, gr3, YPOS2
 586 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 587 => b"01000_0011_01_000000000000", -- mul, gr3
 588 => b"00000_0000_00_000000001111", -- 15
 589 => b"00010_0011_00_001101000100", -- add, gr3, XPOS2
 590 => b"10000_0011_00_000000000000", -- tpoint, gr3
 591 => b"01110_0010_00_000000000000", -- twrite, gr2
 592 => b"00000_0000_01_000000000000", -- load, gr0
 593 => b"00000_0000_00_000000000001", -- 1
 594 => b"00001_0000_10_001100101111", -- store, gr0, P2BOMB1ACTIVE
 595 => b"00001_0011_10_001100101101", -- store, gr3, P2BOMB1POS
 596 => b"00000_0000_01_000000000000", -- load, gr0
 597 => b"00000_0000_00_000000010000", -- 16
 598 => b"00001_0000_10_001100101110", -- store, gr0, P2BOMB1TIME
 599 => b"00100_0000_01_000000000000", -- jump
 600 => b"00000_0000_00_001001000001", -- P2INCREASEBOMBCOUNTER
 601 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 602 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 603 => b"00000_0011_00_001101000101", -- load, gr3, YPOS2
 604 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 605 => b"01000_0011_01_000000000000", -- mul, gr3
 606 => b"00000_0000_00_000000001111", -- 15
 607 => b"00010_0011_00_001101000100", -- add, gr3, XPOS2
 608 => b"10000_0011_00_000000000000", -- tpoint, gr3
 609 => b"01110_0010_00_000000000000", -- twrite, gr2
 610 => b"00000_0000_01_000000000000", -- load, gr0
 611 => b"00000_0000_00_000000000001", -- 1
 612 => b"00001_0000_10_001100110101", -- store, gr0, P2BOMB2ACTIVE
 613 => b"00001_0011_10_001100110011", -- store, gr3, P2BOMB2POS
 614 => b"00000_0000_01_000000000000", -- load, gr0
 615 => b"00000_0000_00_000000010000", -- 16
 616 => b"00001_0000_10_001100110100", -- store, gr0, P2BOMB2TIME
 617 => b"00100_0000_01_000000000000", -- jump
 618 => b"00000_0000_00_001001000001", -- P2INCREASEBOMBCOUNTER
 619 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 620 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 621 => b"00000_0011_00_001101000101", -- load, gr3, YPOS2
 622 => b"00000_0010_00_001101001101", -- load, gr2, EGG
 623 => b"01000_0011_01_000000000000", -- mul, gr3
 624 => b"00000_0000_00_000000001111", -- 15
 625 => b"00010_0011_00_001101000100", -- add, gr3, XPOS2
 626 => b"10000_0011_00_000000000000", -- tpoint, gr3
 627 => b"01110_0010_00_000000000000", -- twrite, gr2
 628 => b"00000_0000_01_000000000000", -- load, gr0
 629 => b"00000_0000_00_000000000001", -- 1
 630 => b"00001_0000_10_001100111011", -- store, gr0, P2BOMB3ACTIVE
 631 => b"00001_0011_10_001100111001", -- store, gr3, P2BOMB3POS
 632 => b"00000_0000_01_000000000000", -- load, gr0
 633 => b"00000_0000_00_000000010000", -- 16
 634 => b"00001_0000_10_001100111010", -- store, gr0, P2BOMB3TIME
 635 => b"00100_0000_01_000000000000", -- jump
 636 => b"00000_0000_00_001001000001", -- P2INCREASEBOMBCOUNTER
 637 => b"00100_0000_01_000000000000", -- jump
 638 => b"00000_0000_00_001100011001", -- COUNT1
 639 => b"10001_0000_01_000000000000", -- joy1r
 640 => b"00000_0000_00_001010010001", -- P1R
 641 => b"10011_0000_01_000000000000", -- joy1l
 642 => b"00000_0000_00_001010110011", -- P1L
 643 => b"10010_0000_01_000000000000", -- joy1u
 644 => b"00000_0000_00_001010100010", -- P1U
 645 => b"10100_0000_01_000000000000", -- joy1d
 646 => b"00000_0000_00_001011000100", -- P1D
 647 => b"10110_0000_01_000000000000", -- joy2r
 648 => b"00000_0000_00_001011010101", -- P2R
 649 => b"11000_0000_01_000000000000", -- joy2l
 650 => b"00000_0000_00_001011110111", -- P2L
 651 => b"10111_0000_01_000000000000", -- joy2u
 652 => b"00000_0000_00_001011100110", -- P2U
 653 => b"11001_0000_01_000000000000", -- joy2d
 654 => b"00000_0000_00_001100001000", -- P2D
 655 => b"00100_0000_01_000000000000", -- jump
 656 => b"00000_0000_00_000000000010", -- CONTROL_R
 657 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 658 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 659 => b"00000_0000_00_001101000011", -- load, gr0, YPOS1
 660 => b"01000_0000_01_000000000000", -- mul, gr0
 661 => b"00000_0000_00_000000001111", -- 15
 662 => b"00010_0000_00_001101000010", -- add, gr0, XPOS1
 663 => b"00010_0000_01_000000000000", -- add, gr0
 664 => b"00000_0000_00_000000000001", -- 1
 665 => b"10000_0000_00_000000000000", -- tpoint, gr0
 666 => b"01111_0001_00_000000000000", -- tread, gr1
 667 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 668 => b"00111_0000_01_000000000000", -- bne
 669 => b"00000_0000_00_001010000011", -- J1
 670 => b"00010_1100_01_000000000000", -- add, gr12
 671 => b"00000_0000_00_000000000001", -- 1
 672 => b"00100_0000_01_000000000000", -- jump
 673 => b"00000_0000_00_001010000011", -- J1
 674 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 675 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 676 => b"00000_0000_00_001101000011", -- load, gr0, YPOS1
 677 => b"00011_0000_01_000000000000", -- sub, gr0
 678 => b"00000_0000_00_000000000001", -- 1
 679 => b"01000_0000_01_000000000000", -- mul, gr0
 680 => b"00000_0000_00_000000001111", -- 15
 681 => b"00010_0000_00_001101000010", -- add, gr0, XPOS1
 682 => b"10000_0000_00_000000000000", -- tpoint, gr0
 683 => b"01111_0001_00_000000000000", -- tread, gr1
 684 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 685 => b"00111_0000_01_000000000000", -- bne
 686 => b"00000_0000_00_001010000111", -- J2
 687 => b"00011_1101_01_000000000000", -- sub, gr13
 688 => b"00000_0000_00_000000000001", -- 1
 689 => b"00100_0000_01_000000000000", -- jump
 690 => b"00000_0000_00_001010000111", -- J2
 691 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 692 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 693 => b"00000_0000_00_001101000011", -- load, gr0, YPOS1
 694 => b"01000_0000_01_000000000000", -- mul, gr0
 695 => b"00000_0000_00_000000001111", -- 15
 696 => b"00010_0000_00_001101000010", -- add, gr0, XPOS1
 697 => b"00011_0000_01_000000000000", -- sub, gr0
 698 => b"00000_0000_00_000000000001", -- 1
 699 => b"10000_0000_00_000000000000", -- tpoint, gr0
 700 => b"01111_0001_00_000000000000", -- tread, gr1
 701 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 702 => b"00111_0000_01_000000000000", -- bne
 703 => b"00000_0000_00_001010000011", -- J1
 704 => b"00011_1100_01_000000000000", -- sub, gr12
 705 => b"00000_0000_00_000000000001", -- 1
 706 => b"00100_0000_01_000000000000", -- jump
 707 => b"00000_0000_00_001010000011", -- J1
 708 => b"00001_1100_10_001101000010", -- store, gr12, XPOS1
 709 => b"00001_1101_10_001101000011", -- store, gr13, YPOS1
 710 => b"00000_0000_00_001101000011", -- load, gr0, YPOS1
 711 => b"00010_0000_01_000000000000", -- add, gr0
 712 => b"00000_0000_00_000000000001", -- 1
 713 => b"01000_0000_01_000000000000", -- mul, gr0
 714 => b"00000_0000_00_000000001111", -- 15
 715 => b"00010_0000_00_001101000010", -- add, gr0, XPOS1
 716 => b"10000_0000_00_000000000000", -- tpoint, gr0
 717 => b"01111_0001_00_000000000000", -- tread, gr1
 718 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 719 => b"00111_0000_01_000000000000", -- bne
 720 => b"00000_0000_00_001010000111", -- J2
 721 => b"00010_1101_01_000000000000", -- add, gr13
 722 => b"00000_0000_00_000000000001", -- 1
 723 => b"00100_0000_01_000000000000", -- jump
 724 => b"00000_0000_00_001010000111", -- J2
 725 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 726 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 727 => b"00000_0000_00_001101000101", -- load, gr0, YPOS2
 728 => b"01000_0000_01_000000000000", -- mul, gr0
 729 => b"00000_0000_00_000000001111", -- 15
 730 => b"00010_0000_00_001101000100", -- add, gr0, XPOS2
 731 => b"00010_0000_01_000000000000", -- add, gr0
 732 => b"00000_0000_00_000000000001", -- 1
 733 => b"10000_0000_00_000000000000", -- tpoint, gr0
 734 => b"01111_0001_00_000000000000", -- tread, gr1
 735 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 736 => b"00111_0000_01_000000000000", -- bne
 737 => b"00000_0000_00_001010001011", -- J3
 738 => b"00010_1110_01_000000000000", -- add, gr14
 739 => b"00000_0000_00_000000000001", -- 1
 740 => b"00100_0000_01_000000000000", -- jump
 741 => b"00000_0000_00_001010001011", -- J3
 742 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 743 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 744 => b"00000_0000_00_001101000101", -- load, gr0, YPOS2
 745 => b"00011_0000_01_000000000000", -- sub, gr0
 746 => b"00000_0000_00_000000000001", -- 1
 747 => b"01000_0000_01_000000000000", -- mul, gr0
 748 => b"00000_0000_00_000000001111", -- 15
 749 => b"00010_0000_00_001101000100", -- add, gr0, XPOS2
 750 => b"10000_0000_00_000000000000", -- tpoint, gr0
 751 => b"01111_0001_00_000000000000", -- tread, gr1
 752 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 753 => b"00111_0000_01_000000000000", -- bne
 754 => b"00000_0000_00_000000000010", -- CONTROL_R
 755 => b"00011_1111_01_000000000000", -- sub, gr15
 756 => b"00000_0000_00_000000000001", -- 1
 757 => b"00100_0000_01_000000000000", -- jump
 758 => b"00000_0000_00_000000000010", -- CONTROL_R
 759 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 760 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 761 => b"00000_0000_00_001101000101", -- load, gr0, YPOS2
 762 => b"01000_0000_01_000000000000", -- mul, gr0
 763 => b"00000_0000_00_000000001111", -- 15
 764 => b"00010_0000_00_001101000100", -- add, gr0, XPOS2
 765 => b"00011_0000_01_000000000000", -- sub, gr0
 766 => b"00000_0000_00_000000000001", -- 1
 767 => b"10000_0000_00_000000000000", -- tpoint, gr0
 768 => b"01111_0001_00_000000000000", -- tread, gr1
 769 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 770 => b"00111_0000_01_000000000000", -- bne
 771 => b"00000_0000_00_001010001011", -- J3
 772 => b"00011_1110_01_000000000000", -- sub, gr14
 773 => b"00000_0000_00_000000000001", -- 1
 774 => b"00100_0000_01_000000000000", -- jump
 775 => b"00000_0000_00_001010001011", -- J3
 776 => b"00001_1110_10_001101000100", -- store, gr14, XPOS2
 777 => b"00001_1111_10_001101000101", -- store, gr15, YPOS2
 778 => b"00000_0000_00_001101000101", -- load, gr0, YPOS2
 779 => b"00010_0000_01_000000000000", -- add, gr0
 780 => b"00000_0000_00_000000000001", -- 1
 781 => b"01000_0000_01_000000000000", -- mul, gr0
 782 => b"00000_0000_00_000000001111", -- 15
 783 => b"00010_0000_00_001101000100", -- add, gr0, XPOS2
 784 => b"10000_0000_00_000000000000", -- tpoint, gr0
 785 => b"01111_0001_00_000000000000", -- tread, gr1
 786 => b"00011_0001_00_001101001001", -- sub, gr1, GRASS
 787 => b"00111_0000_01_000000000000", -- bne
 788 => b"00000_0000_00_000000000010", -- CONTROL_R
 789 => b"00010_1111_01_000000000000", -- add, gr15
 790 => b"00000_0000_00_000000000001", -- 1
 791 => b"00100_0000_01_000000000000", -- jump
 792 => b"00000_0000_00_000000000010", -- CONTROL_R
 793 => b"00100_0000_01_000000000000", -- jump
 794 => b"00000_0000_00_001001111111", -- COUNT_R
 795 => b"00000_0000_00_000000000000", -- 0
 796 => b"00000_0000_00_000000000000", -- 0
 797 => b"00000_0000_00_000000000000", -- 0
 798 => b"00000_0000_00_000000000000", -- 0
 799 => b"00000_0000_00_000000000000", -- 0
 800 => b"00000_0000_00_000000000000", -- 0
 801 => b"00000_0000_00_000000000000", -- 0
 802 => b"00000_0000_00_000000000000", -- 0
 803 => b"00000_0000_00_000000000000", -- 0
 804 => b"00000_0000_00_000000000000", -- 0
 805 => b"00000_0000_00_000000000000", -- 0
 806 => b"00000_0000_00_000000000000", -- 0
 807 => b"00000_0000_00_000000000000", -- 0
 808 => b"00000_0000_00_000000000000", -- 0
 809 => b"00000_0000_00_000000000000", -- 0
 810 => b"00000_0000_00_000000000000", -- 0
 811 => b"00000_0000_00_000000000000", -- 0
 812 => b"00000_0000_00_000000000000", -- 0
 813 => b"00000_0000_00_000000000000", -- 0
 814 => b"00000_0000_00_000000000000", -- 0
 815 => b"00000_0000_00_000000000000", -- 0
 816 => b"00000_0000_00_000000000000", -- 0
 817 => b"00000_0000_00_000000000000", -- 0
 818 => b"00000_0000_00_000000000000", -- 0
 819 => b"00000_0000_00_000000000000", -- 0
 820 => b"00000_0000_00_000000000000", -- 0
 821 => b"00000_0000_00_000000000000", -- 0
 822 => b"00000_0000_00_000000000000", -- 0
 823 => b"00000_0000_00_000000000000", -- 0
 824 => b"00000_0000_00_000000000000", -- 0
 825 => b"00000_0000_00_000000000000", -- 0
 826 => b"00000_0000_00_000000000000", -- 0
 827 => b"00000_0000_00_000000000000", -- 0
 828 => b"00000_0000_00_000000000000", -- 0
 829 => b"00000_0000_00_000000000000", -- 0
 830 => b"00000_0000_00_000000000000", -- 0
 831 => b"00000_0000_00_000000000000", -- 0
 832 => b"00000_0000_00_000000000000", -- 0
 833 => b"00000_0000_00_000000000011", -- 3
 834 => b"00000_0000_00_000000000000", -- 0
 835 => b"00000_0000_00_000000000000", -- 0
 836 => b"00000_0000_00_000000000000", -- 0
 837 => b"00000_0000_00_000000000000", -- 0
 838 => b"00000_0000_00_000000000000", -- 0
 839 => b"00000_0000_00_000000000000", -- 0
 840 => b"00000_0000_00_000000000000", -- 0
 841 => b"00000_0000_00_000000000000", -- 0
 842 => b"00000_0000_00_000000000001", -- 1
 843 => b"00000_0000_00_000000000010", -- 2
 844 => b"00000_0000_00_000000000011", -- 3
 845 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
