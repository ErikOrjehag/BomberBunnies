library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr
0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000000100101", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000000001000", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000000010", -- MAIN
   8 => b"10101_0000_01_000000000000", -- btn1
   9 => b"00000_0000_00_000000001110", -- BTN1
  10 => b"11010_0000_01_000000000000", -- btn2
  11 => b"00000_0000_00_000000011001", -- BTN2
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000000000110", -- BUTTON_R
  14 => b"00001_1100_10_000011001000", -- store, gr12, XPOS1
  15 => b"00001_1101_10_000011001001", -- store, gr13, YPOS1
  16 => b"00000_0011_00_000011001001", -- load, gr3, YPOS1
  17 => b"00000_0010_00_000011000111", -- load, gr2, EGG
  18 => b"01000_0011_01_000000000000", -- mul, gr3
  19 => b"00000_0000_00_000000001111", -- 15
  20 => b"00010_0011_00_000011001000", -- add, gr3, XPOS1
  21 => b"10000_0011_00_000000000000", -- tpoint, gr3
  22 => b"01110_0010_00_000000000000", -- twrite, gr2
  23 => b"00100_0000_01_000000000000", -- jump
  24 => b"00000_0000_00_000000001010", -- BTN1_R
  25 => b"00001_1110_10_000011001010", -- store, gr14, XPOS2
  26 => b"00001_1111_10_000011001011", -- store, gr15, YPOS2
  27 => b"00000_0011_00_000011001011", -- load, gr3, YPOS2
  28 => b"00000_0010_00_000011000111", -- load, gr2, EGG
  29 => b"01000_0011_01_000000000000", -- mul, gr3
  30 => b"00000_0000_00_000000001111", -- 15
  31 => b"00010_0011_00_000011001010", -- add, gr3, XPOS2
  32 => b"10000_0011_00_000000000000", -- tpoint, gr3
  33 => b"01110_0010_00_000000000000", -- twrite, gr2
  34 => b"00100_0000_01_000000000000", -- jump
  35 => b"00000_0000_00_000000001100", -- BTN2_R
  36 => b"00000_0000_00_000000000000", -- 0
  37 => b"00100_0000_01_000000000000", -- jump
  38 => b"00000_0000_00_000011000001", -- COUNT1
  39 => b"10001_0000_01_000000000000", -- joy1r
  40 => b"00000_0000_00_000000111001", -- P1R
  41 => b"10011_0000_01_000000000000", -- joy1l
  42 => b"00000_0000_00_000001011011", -- P1L
  43 => b"10010_0000_01_000000000000", -- joy1u
  44 => b"00000_0000_00_000001001010", -- P1U
  45 => b"10100_0000_01_000000000000", -- joy1d
  46 => b"00000_0000_00_000001101100", -- P1D
  47 => b"10110_0000_01_000000000000", -- joy2r
  48 => b"00000_0000_00_000001111101", -- P2R
  49 => b"11000_0000_01_000000000000", -- joy2l
  50 => b"00000_0000_00_000010011111", -- P2L
  51 => b"10111_0000_01_000000000000", -- joy2u
  52 => b"00000_0000_00_000010001110", -- P2U
  53 => b"11001_0000_01_000000000000", -- joy2d
  54 => b"00000_0000_00_000010110000", -- P2D
  55 => b"00100_0000_01_000000000000", -- jump
  56 => b"00000_0000_00_000000000100", -- CONTROL_R
  57 => b"00001_1100_10_000011001000", -- store, gr12, XPOS1
  58 => b"00001_1101_10_000011001001", -- store, gr13, YPOS1
  59 => b"00000_0000_00_000011001001", -- load, gr0, YPOS1
  60 => b"01000_0000_01_000000000000", -- mul, gr0
  61 => b"00000_0000_00_000000001111", -- 15
  62 => b"00010_0000_00_000011001000", -- add, gr0, XPOS1
  63 => b"00010_0000_01_000000000000", -- add, gr0
  64 => b"00000_0000_00_000000000001", -- 1
  65 => b"10000_0000_00_000000000000", -- tpoint, gr0
  66 => b"01111_0001_00_000000000000", -- tread, gr1
  67 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
  68 => b"00111_0000_01_000000000000", -- bne
  69 => b"00000_0000_00_000000101011", -- J1
  70 => b"00010_1100_01_000000000000", -- add, gr12
  71 => b"00000_0000_00_000000000001", -- 1
  72 => b"00100_0000_01_000000000000", -- jump
  73 => b"00000_0000_00_000000101011", -- J1
  74 => b"00001_1100_10_000011001000", -- store, gr12, XPOS1
  75 => b"00001_1101_10_000011001001", -- store, gr13, YPOS1
  76 => b"00000_0000_00_000011001001", -- load, gr0, YPOS1
  77 => b"00011_0000_01_000000000000", -- sub, gr0
  78 => b"00000_0000_00_000000000001", -- 1
  79 => b"01000_0000_01_000000000000", -- mul, gr0
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"00010_0000_00_000011001000", -- add, gr0, XPOS1
  82 => b"10000_0000_00_000000000000", -- tpoint, gr0
  83 => b"01111_0001_00_000000000000", -- tread, gr1
  84 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
  85 => b"00111_0000_01_000000000000", -- bne
  86 => b"00000_0000_00_000000101111", -- J2
  87 => b"00011_1101_01_000000000000", -- sub, gr13
  88 => b"00000_0000_00_000000000001", -- 1
  89 => b"00100_0000_01_000000000000", -- jump
  90 => b"00000_0000_00_000000101111", -- J2
  91 => b"00001_1100_10_000011001000", -- store, gr12, XPOS1
  92 => b"00001_1101_10_000011001001", -- store, gr13, YPOS1
  93 => b"00000_0000_00_000011001001", -- load, gr0, YPOS1
  94 => b"01000_0000_01_000000000000", -- mul, gr0
  95 => b"00000_0000_00_000000001111", -- 15
  96 => b"00010_0000_00_000011001000", -- add, gr0, XPOS1
  97 => b"00011_0000_01_000000000000", -- sub, gr0
  98 => b"00000_0000_00_000000000001", -- 1
  99 => b"10000_0000_00_000000000000", -- tpoint, gr0
 100 => b"01111_0001_00_000000000000", -- tread, gr1
 101 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 102 => b"00111_0000_01_000000000000", -- bne
 103 => b"00000_0000_00_000000101011", -- J1
 104 => b"00011_1100_01_000000000000", -- sub, gr12
 105 => b"00000_0000_00_000000000001", -- 1
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000000101011", -- J1
 108 => b"00001_1100_10_000011001000", -- store, gr12, XPOS1
 109 => b"00001_1101_10_000011001001", -- store, gr13, YPOS1
 110 => b"00000_0000_00_000011001001", -- load, gr0, YPOS1
 111 => b"00010_0000_01_000000000000", -- add, gr0
 112 => b"00000_0000_00_000000000001", -- 1
 113 => b"01000_0000_01_000000000000", -- mul, gr0
 114 => b"00000_0000_00_000000001111", -- 15
 115 => b"00010_0000_00_000011001000", -- add, gr0, XPOS1
 116 => b"10000_0000_00_000000000000", -- tpoint, gr0
 117 => b"01111_0001_00_000000000000", -- tread, gr1
 118 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 119 => b"00111_0000_01_000000000000", -- bne
 120 => b"00000_0000_00_000000101111", -- J2
 121 => b"00010_1101_01_000000000000", -- add, gr13
 122 => b"00000_0000_00_000000000001", -- 1
 123 => b"00100_0000_01_000000000000", -- jump
 124 => b"00000_0000_00_000000101111", -- J2
 125 => b"00001_1110_10_000011001010", -- store, gr14, XPOS2
 126 => b"00001_1111_10_000011001011", -- store, gr15, YPOS2
 127 => b"00000_0000_00_000011001011", -- load, gr0, YPOS2
 128 => b"01000_0000_01_000000000000", -- mul, gr0
 129 => b"00000_0000_00_000000001111", -- 15
 130 => b"00010_0000_00_000011001010", -- add, gr0, XPOS2
 131 => b"00010_0000_01_000000000000", -- add, gr0
 132 => b"00000_0000_00_000000000001", -- 1
 133 => b"10000_0000_00_000000000000", -- tpoint, gr0
 134 => b"01111_0001_00_000000000000", -- tread, gr1
 135 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 136 => b"00111_0000_01_000000000000", -- bne
 137 => b"00000_0000_00_000000110011", -- J3
 138 => b"00010_1110_01_000000000000", -- add, gr14
 139 => b"00000_0000_00_000000000001", -- 1
 140 => b"00100_0000_01_000000000000", -- jump
 141 => b"00000_0000_00_000000110011", -- J3
 142 => b"00001_1110_10_000011001010", -- store, gr14, XPOS2
 143 => b"00001_1111_10_000011001011", -- store, gr15, YPOS2
 144 => b"00000_0000_00_000011001011", -- load, gr0, YPOS2
 145 => b"00011_0000_01_000000000000", -- sub, gr0
 146 => b"00000_0000_00_000000000001", -- 1
 147 => b"01000_0000_01_000000000000", -- mul, gr0
 148 => b"00000_0000_00_000000001111", -- 15
 149 => b"00010_0000_00_000011001010", -- add, gr0, XPOS2
 150 => b"10000_0000_00_000000000000", -- tpoint, gr0
 151 => b"01111_0001_00_000000000000", -- tread, gr1
 152 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 153 => b"00111_0000_01_000000000000", -- bne
 154 => b"00000_0000_00_000000000100", -- CONTROL_R
 155 => b"00011_1111_01_000000000000", -- sub, gr15
 156 => b"00000_0000_00_000000000001", -- 1
 157 => b"00100_0000_01_000000000000", -- jump
 158 => b"00000_0000_00_000000000100", -- CONTROL_R
 159 => b"00001_1110_10_000011001010", -- store, gr14, XPOS2
 160 => b"00001_1111_10_000011001011", -- store, gr15, YPOS2
 161 => b"00000_0000_00_000011001011", -- load, gr0, YPOS2
 162 => b"01000_0000_01_000000000000", -- mul, gr0
 163 => b"00000_0000_00_000000001111", -- 15
 164 => b"00010_0000_00_000011001010", -- add, gr0, XPOS2
 165 => b"00011_0000_01_000000000000", -- sub, gr0
 166 => b"00000_0000_00_000000000001", -- 1
 167 => b"10000_0000_00_000000000000", -- tpoint, gr0
 168 => b"01111_0001_00_000000000000", -- tread, gr1
 169 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 170 => b"00111_0000_01_000000000000", -- bne
 171 => b"00000_0000_00_000000110011", -- J3
 172 => b"00011_1110_01_000000000000", -- sub, gr14
 173 => b"00000_0000_00_000000000001", -- 1
 174 => b"00100_0000_01_000000000000", -- jump
 175 => b"00000_0000_00_000000110011", -- J3
 176 => b"00001_1110_10_000011001010", -- store, gr14, XPOS2
 177 => b"00001_1111_10_000011001011", -- store, gr15, YPOS2
 178 => b"00000_0000_00_000011001011", -- load, gr0, YPOS2
 179 => b"00010_0000_01_000000000000", -- add, gr0
 180 => b"00000_0000_00_000000000001", -- 1
 181 => b"01000_0000_01_000000000000", -- mul, gr0
 182 => b"00000_0000_00_000000001111", -- 15
 183 => b"00010_0000_00_000011001010", -- add, gr0, XPOS2
 184 => b"10000_0000_00_000000000000", -- tpoint, gr0
 185 => b"01111_0001_00_000000000000", -- tread, gr1
 186 => b"00011_0001_00_000011000011", -- sub, gr1, GRASS
 187 => b"00111_0000_01_000000000000", -- bne
 188 => b"00000_0000_00_000000000100", -- CONTROL_R
 189 => b"00010_1111_01_000000000000", -- add, gr15
 190 => b"00000_0000_00_000000000001", -- 1
 191 => b"00100_0000_01_000000000000", -- jump
 192 => b"00000_0000_00_000000000100", -- CONTROL_R
 193 => b"00100_0000_01_000000000000", -- jump
 194 => b"00000_0000_00_000000100111", -- COUNT_R
 195 => b"00000_0000_00_000000000000", -- 0
 196 => b"00000_0000_00_000000000001", -- 1
 197 => b"00000_0000_00_000000000010", -- 2
 198 => b"00000_0000_00_000000000011", -- 3
 199 => b"00000_0000_00_000000000100", -- 4
 200 => b"00000_0000_00_000000000000", -- 0
 201 => b"00000_0000_00_000000000000", -- 0
 202 => b"00000_0000_00_000000000000", -- 0
 203 => b"00000_0000_00_000000000000", -- 0
 204 => b"00000_0000_00_000000000000", -- 0
 205 => b"00000_0000_00_000000000000", -- 0
 206 => b"00000_0000_00_000000000000", -- 0


   


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


