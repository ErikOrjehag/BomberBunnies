library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr




    

0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000010110001", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000001100111", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKBOMBS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000010", -- MAIN
  10 => b"00000_0000_00_000101010001", -- load, gr0, P1BOMBACTIVE
  11 => b"00011_0000_01_000000000000", -- sub, gr0
  12 => b"00000_0000_00_000000000001", -- 1
  13 => b"00111_0000_01_000000000000", -- bne
  14 => b"00000_0000_00_000001100101", -- TICK2
  15 => b"00000_0000_00_000101010000", -- load, gr0, P1BOMBTIME
  16 => b"00011_0000_01_000000000000", -- sub, gr0
  17 => b"00000_0000_00_000000000001", -- 1
  18 => b"00001_0000_10_000101010000", -- store, gr0, P1BOMBTIME
  19 => b"00000_0000_01_000000000000", -- load, gr0
  20 => b"00000_0000_00_000000000000", -- 0
  21 => b"00011_0000_00_000101010000", -- sub, gr0, P1BOMBTIME
  22 => b"00110_0000_01_000000000000", -- beq
  23 => b"00000_0000_00_000000011010", -- EXPLODE1
  24 => b"00100_0000_01_000000000000", -- jump
  25 => b"00000_0000_00_000001100101", -- TICK2
  26 => b"00000_0000_00_000101010101", -- load, gr0, BOMBS1
  27 => b"00011_0000_01_000000000000", -- sub, gr0
  28 => b"00000_0000_00_000000000001", -- 1
  29 => b"00001_0000_10_000101010101", -- store, gr0, BOMBS1
  30 => b"00000_0010_00_000101001111", -- load, gr2, P1BOMBPOS
  31 => b"00000_0011_00_000101011011", -- load, gr3, EXPLOSION
  32 => b"10000_0010_00_000000000000", -- tpoint, gr2
  33 => b"01110_0011_00_000000000000", -- twrite, gr3
  34 => b"00010_0010_01_000000000000", -- add, gr2
  35 => b"00000_0000_00_000000000001", -- 1
  36 => b"10000_0010_00_000000000000", -- tpoint, gr2
  37 => b"01111_0000_00_000000000000", -- tread, gr0
  38 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  39 => b"00110_0000_01_000000000000", -- beq
  40 => b"00000_0000_00_000000110010", -- P1LEFT
  41 => b"01110_0011_00_000000000000", -- twrite, gr3
  42 => b"00010_0010_01_000000000000", -- add, gr2
  43 => b"00000_0000_00_000000000001", -- 1
  44 => b"10000_0010_00_000000000000", -- tpoint, gr2
  45 => b"01111_0000_00_000000000000", -- tread, gr0
  46 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  47 => b"00110_0000_01_000000000000", -- beq
  48 => b"00000_0000_00_000000110010", -- P1LEFT
  49 => b"01110_0011_00_000000000000", -- twrite, gr3
  50 => b"00000_0010_00_000101001111", -- load, gr2, P1BOMBPOS
  51 => b"00011_0010_01_000000000000", -- sub, gr2
  52 => b"00000_0000_00_000000000001", -- 1
  53 => b"10000_0010_00_000000000000", -- tpoint, gr2
  54 => b"01111_0000_00_000000000000", -- tread, gr0
  55 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  56 => b"00110_0000_01_000000000000", -- beq
  57 => b"00000_0000_00_000001000011", -- P1DOWN
  58 => b"01110_0011_00_000000000000", -- twrite, gr3
  59 => b"00011_0010_01_000000000000", -- sub, gr2
  60 => b"00000_0000_00_000000000001", -- 1
  61 => b"10000_0010_00_000000000000", -- tpoint, gr2
  62 => b"01111_0000_00_000000000000", -- tread, gr0
  63 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  64 => b"00110_0000_01_000000000000", -- beq
  65 => b"00000_0000_00_000001000011", -- P1DOWN
  66 => b"01110_0011_00_000000000000", -- twrite, gr3
  67 => b"00000_0010_00_000101001111", -- load, gr2, P1BOMBPOS
  68 => b"00010_0010_01_000000000000", -- add, gr2
  69 => b"00000_0000_00_000000001111", -- 15
  70 => b"10000_0010_00_000000000000", -- tpoint, gr2
  71 => b"01111_0000_00_000000000000", -- tread, gr0
  72 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  73 => b"00110_0000_01_000000000000", -- beq
  74 => b"00000_0000_00_000001010100", -- P1UP
  75 => b"01110_0011_00_000000000000", -- twrite, gr3
  76 => b"00010_0010_01_000000000000", -- add, gr2
  77 => b"00000_0000_00_000000001111", -- 15
  78 => b"10000_0010_00_000000000000", -- tpoint, gr2
  79 => b"01111_0000_00_000000000000", -- tread, gr0
  80 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  81 => b"00110_0000_01_000000000000", -- beq
  82 => b"00000_0000_00_000001010100", -- P1UP
  83 => b"01110_0011_00_000000000000", -- twrite, gr3
  84 => b"00000_0010_00_000101001111", -- load, gr2, P1BOMBPOS
  85 => b"00011_0010_01_000000000000", -- sub, gr2
  86 => b"00000_0000_00_000000001111", -- 15
  87 => b"10000_0010_00_000000000000", -- tpoint, gr2
  88 => b"01111_0000_00_000000000000", -- tread, gr0
  89 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  90 => b"00110_0000_01_000000000000", -- beq
  91 => b"00000_0000_00_000001100101", -- TICK2
  92 => b"01110_0011_00_000000000000", -- twrite, gr3
  93 => b"00011_0010_01_000000000000", -- sub, gr2
  94 => b"00000_0000_00_000000001111", -- 15
  95 => b"10000_0010_00_000000000000", -- tpoint, gr2
  96 => b"01111_0000_00_000000000000", -- tread, gr0
  97 => b"00011_0000_00_000101011001", -- sub, gr0, WALL
  98 => b"00110_0000_01_000000000000", -- beq
  99 => b"00000_0000_00_000001100101", -- TICK2
 100 => b"01110_0011_00_000000000000", -- twrite, gr3
 101 => b"00100_0000_01_000000000000", -- jump
 102 => b"00000_0000_00_000000001000", -- TICKBOMBS_R
 103 => b"10101_0000_01_000000000000", -- btn1
 104 => b"00000_0000_00_000001101101", -- BTN1
 105 => b"11010_0000_01_000000000000", -- btn2
 106 => b"00000_0000_00_000010010010", -- BTN2
 107 => b"00100_0000_01_000000000000", -- jump
 108 => b"00000_0000_00_000000000110", -- BUTTON_R
 109 => b"00000_0000_00_000101010101", -- load, gr0, BOMBS1
 110 => b"00011_0000_00_000101010111", -- sub, gr0, MAXBOMBS
 111 => b"00110_0000_01_000000000000", -- beq
 112 => b"00000_0000_00_000001101001", -- BTN1_R
 113 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 114 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 115 => b"00000_0000_00_000101011110", -- load, gr0, YPOS1
 116 => b"01000_0000_01_000000000000", -- mul, gr0
 117 => b"00000_0000_00_000000001111", -- 15
 118 => b"00010_0000_00_000101011101", -- add, gr0, XPOS1
 119 => b"10000_0000_00_000000000000", -- tpoint, gr0
 120 => b"01111_0001_00_000000000000", -- tread, gr1
 121 => b"00011_0001_00_000101011100", -- sub, gr1, EGG
 122 => b"00110_0000_01_000000000000", -- beq
 123 => b"00000_0000_00_000001101011", -- BTN2_R
 124 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 125 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 126 => b"00000_0011_00_000101011110", -- load, gr3, YPOS1
 127 => b"00000_0010_00_000101011100", -- load, gr2, EGG
 128 => b"01000_0011_01_000000000000", -- mul, gr3
 129 => b"00000_0000_00_000000001111", -- 15
 130 => b"00010_0011_00_000101011101", -- add, gr3, XPOS1
 131 => b"10000_0011_00_000000000000", -- tpoint, gr3
 132 => b"01110_0010_00_000000000000", -- twrite, gr2
 133 => b"00000_0000_01_000000000000", -- load, gr0
 134 => b"00000_0000_00_000000000001", -- 1
 135 => b"00001_0000_10_000101010001", -- store, gr0, P1BOMBACTIVE
 136 => b"00001_0011_10_000101001111", -- store, gr3, P1BOMBPOS
 137 => b"00000_0000_01_000000000000", -- load, gr0
 138 => b"00000_0000_00_000000010000", -- 16
 139 => b"00001_0000_10_000101010000", -- store, gr0, P1BOMBTIME
 140 => b"00000_0000_00_000101010101", -- load, gr0, BOMBS1
 141 => b"00010_0000_01_000000000000", -- add, gr0
 142 => b"00000_0000_00_000000000001", -- 1
 143 => b"00001_0000_10_000101010101", -- store, gr0, BOMBS1
 144 => b"00100_0000_01_000000000000", -- jump
 145 => b"00000_0000_00_000001101001", -- BTN1_R
 146 => b"00000_0000_00_000101010110", -- load, gr0, BOMBS2
 147 => b"00011_0000_00_000101010111", -- sub, gr0, MAXBOMBS
 148 => b"00110_0000_01_000000000000", -- beq
 149 => b"00000_0000_00_000001101011", -- BTN2_R
 150 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 151 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 152 => b"00000_0000_00_000101100000", -- load, gr0, YPOS2
 153 => b"01000_0000_01_000000000000", -- mul, gr0
 154 => b"00000_0000_00_000000001111", -- 15
 155 => b"00010_0000_00_000101011111", -- add, gr0, XPOS2
 156 => b"10000_0000_00_000000000000", -- tpoint, gr0
 157 => b"01111_0001_00_000000000000", -- tread, gr1
 158 => b"00011_0001_00_000101011100", -- sub, gr1, EGG
 159 => b"00110_0000_01_000000000000", -- beq
 160 => b"00000_0000_00_000001101011", -- BTN2_R
 161 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 162 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 163 => b"00000_0011_00_000101100000", -- load, gr3, YPOS2
 164 => b"00000_0010_00_000101011100", -- load, gr2, EGG
 165 => b"01000_0011_01_000000000000", -- mul, gr3
 166 => b"00000_0000_00_000000001111", -- 15
 167 => b"00010_0011_00_000101011111", -- add, gr3, XPOS2
 168 => b"10000_0011_00_000000000000", -- tpoint, gr3
 169 => b"01110_0010_00_000000000000", -- twrite, gr2
 170 => b"00000_0000_00_000101010110", -- load, gr0, BOMBS2
 171 => b"00010_0000_01_000000000000", -- add, gr0
 172 => b"00000_0000_00_000000000001", -- 1
 173 => b"00001_0000_10_000101010110", -- store, gr0, BOMBS2
 174 => b"00100_0000_01_000000000000", -- jump
 175 => b"00000_0000_00_000001101011", -- BTN2_R
 176 => b"00000_0000_00_000000000000", -- 0
 177 => b"00100_0000_01_000000000000", -- jump
 178 => b"00000_0000_00_000101001101", -- COUNT1
 179 => b"10001_0000_01_000000000000", -- joy1r
 180 => b"00000_0000_00_000011000101", -- P1R
 181 => b"10011_0000_01_000000000000", -- joy1l
 182 => b"00000_0000_00_000011100111", -- P1L
 183 => b"10010_0000_01_000000000000", -- joy1u
 184 => b"00000_0000_00_000011010110", -- P1U
 185 => b"10100_0000_01_000000000000", -- joy1d
 186 => b"00000_0000_00_000011111000", -- P1D
 187 => b"10110_0000_01_000000000000", -- joy2r
 188 => b"00000_0000_00_000100001001", -- P2R
 189 => b"11000_0000_01_000000000000", -- joy2l
 190 => b"00000_0000_00_000100101011", -- P2L
 191 => b"10111_0000_01_000000000000", -- joy2u
 192 => b"00000_0000_00_000100011010", -- P2U
 193 => b"11001_0000_01_000000000000", -- joy2d
 194 => b"00000_0000_00_000100111100", -- P2D
 195 => b"00100_0000_01_000000000000", -- jump
 196 => b"00000_0000_00_000000000100", -- CONTROL_R
 197 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 198 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 199 => b"00000_0000_00_000101011110", -- load, gr0, YPOS1
 200 => b"01000_0000_01_000000000000", -- mul, gr0
 201 => b"00000_0000_00_000000001111", -- 15
 202 => b"00010_0000_00_000101011101", -- add, gr0, XPOS1
 203 => b"00010_0000_01_000000000000", -- add, gr0
 204 => b"00000_0000_00_000000000001", -- 1
 205 => b"10000_0000_00_000000000000", -- tpoint, gr0
 206 => b"01111_0001_00_000000000000", -- tread, gr1
 207 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 208 => b"00111_0000_01_000000000000", -- bne
 209 => b"00000_0000_00_000010110111", -- J1
 210 => b"00010_1100_01_000000000000", -- add, gr12
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00100_0000_01_000000000000", -- jump
 213 => b"00000_0000_00_000010110111", -- J1
 214 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 215 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 216 => b"00000_0000_00_000101011110", -- load, gr0, YPOS1
 217 => b"00011_0000_01_000000000000", -- sub, gr0
 218 => b"00000_0000_00_000000000001", -- 1
 219 => b"01000_0000_01_000000000000", -- mul, gr0
 220 => b"00000_0000_00_000000001111", -- 15
 221 => b"00010_0000_00_000101011101", -- add, gr0, XPOS1
 222 => b"10000_0000_00_000000000000", -- tpoint, gr0
 223 => b"01111_0001_00_000000000000", -- tread, gr1
 224 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 225 => b"00111_0000_01_000000000000", -- bne
 226 => b"00000_0000_00_000010111011", -- J2
 227 => b"00011_1101_01_000000000000", -- sub, gr13
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00100_0000_01_000000000000", -- jump
 230 => b"00000_0000_00_000010111011", -- J2
 231 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 232 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 233 => b"00000_0000_00_000101011110", -- load, gr0, YPOS1
 234 => b"01000_0000_01_000000000000", -- mul, gr0
 235 => b"00000_0000_00_000000001111", -- 15
 236 => b"00010_0000_00_000101011101", -- add, gr0, XPOS1
 237 => b"00011_0000_01_000000000000", -- sub, gr0
 238 => b"00000_0000_00_000000000001", -- 1
 239 => b"10000_0000_00_000000000000", -- tpoint, gr0
 240 => b"01111_0001_00_000000000000", -- tread, gr1
 241 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 242 => b"00111_0000_01_000000000000", -- bne
 243 => b"00000_0000_00_000010110111", -- J1
 244 => b"00011_1100_01_000000000000", -- sub, gr12
 245 => b"00000_0000_00_000000000001", -- 1
 246 => b"00100_0000_01_000000000000", -- jump
 247 => b"00000_0000_00_000010110111", -- J1
 248 => b"00001_1100_10_000101011101", -- store, gr12, XPOS1
 249 => b"00001_1101_10_000101011110", -- store, gr13, YPOS1
 250 => b"00000_0000_00_000101011110", -- load, gr0, YPOS1
 251 => b"00010_0000_01_000000000000", -- add, gr0
 252 => b"00000_0000_00_000000000001", -- 1
 253 => b"01000_0000_01_000000000000", -- mul, gr0
 254 => b"00000_0000_00_000000001111", -- 15
 255 => b"00010_0000_00_000101011101", -- add, gr0, XPOS1
 256 => b"10000_0000_00_000000000000", -- tpoint, gr0
 257 => b"01111_0001_00_000000000000", -- tread, gr1
 258 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 259 => b"00111_0000_01_000000000000", -- bne
 260 => b"00000_0000_00_000010111011", -- J2
 261 => b"00010_1101_01_000000000000", -- add, gr13
 262 => b"00000_0000_00_000000000001", -- 1
 263 => b"00100_0000_01_000000000000", -- jump
 264 => b"00000_0000_00_000010111011", -- J2
 265 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 266 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 267 => b"00000_0000_00_000101100000", -- load, gr0, YPOS2
 268 => b"01000_0000_01_000000000000", -- mul, gr0
 269 => b"00000_0000_00_000000001111", -- 15
 270 => b"00010_0000_00_000101011111", -- add, gr0, XPOS2
 271 => b"00010_0000_01_000000000000", -- add, gr0
 272 => b"00000_0000_00_000000000001", -- 1
 273 => b"10000_0000_00_000000000000", -- tpoint, gr0
 274 => b"01111_0001_00_000000000000", -- tread, gr1
 275 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 276 => b"00111_0000_01_000000000000", -- bne
 277 => b"00000_0000_00_000010111111", -- J3
 278 => b"00010_1110_01_000000000000", -- add, gr14
 279 => b"00000_0000_00_000000000001", -- 1
 280 => b"00100_0000_01_000000000000", -- jump
 281 => b"00000_0000_00_000010111111", -- J3
 282 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 283 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 284 => b"00000_0000_00_000101100000", -- load, gr0, YPOS2
 285 => b"00011_0000_01_000000000000", -- sub, gr0
 286 => b"00000_0000_00_000000000001", -- 1
 287 => b"01000_0000_01_000000000000", -- mul, gr0
 288 => b"00000_0000_00_000000001111", -- 15
 289 => b"00010_0000_00_000101011111", -- add, gr0, XPOS2
 290 => b"10000_0000_00_000000000000", -- tpoint, gr0
 291 => b"01111_0001_00_000000000000", -- tread, gr1
 292 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 293 => b"00111_0000_01_000000000000", -- bne
 294 => b"00000_0000_00_000000000100", -- CONTROL_R
 295 => b"00011_1111_01_000000000000", -- sub, gr15
 296 => b"00000_0000_00_000000000001", -- 1
 297 => b"00100_0000_01_000000000000", -- jump
 298 => b"00000_0000_00_000000000100", -- CONTROL_R
 299 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 300 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 301 => b"00000_0000_00_000101100000", -- load, gr0, YPOS2
 302 => b"01000_0000_01_000000000000", -- mul, gr0
 303 => b"00000_0000_00_000000001111", -- 15
 304 => b"00010_0000_00_000101011111", -- add, gr0, XPOS2
 305 => b"00011_0000_01_000000000000", -- sub, gr0
 306 => b"00000_0000_00_000000000001", -- 1
 307 => b"10000_0000_00_000000000000", -- tpoint, gr0
 308 => b"01111_0001_00_000000000000", -- tread, gr1
 309 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 310 => b"00111_0000_01_000000000000", -- bne
 311 => b"00000_0000_00_000010111111", -- J3
 312 => b"00011_1110_01_000000000000", -- sub, gr14
 313 => b"00000_0000_00_000000000001", -- 1
 314 => b"00100_0000_01_000000000000", -- jump
 315 => b"00000_0000_00_000010111111", -- J3
 316 => b"00001_1110_10_000101011111", -- store, gr14, XPOS2
 317 => b"00001_1111_10_000101100000", -- store, gr15, YPOS2
 318 => b"00000_0000_00_000101100000", -- load, gr0, YPOS2
 319 => b"00010_0000_01_000000000000", -- add, gr0
 320 => b"00000_0000_00_000000000001", -- 1
 321 => b"01000_0000_01_000000000000", -- mul, gr0
 322 => b"00000_0000_00_000000001111", -- 15
 323 => b"00010_0000_00_000101011111", -- add, gr0, XPOS2
 324 => b"10000_0000_00_000000000000", -- tpoint, gr0
 325 => b"01111_0001_00_000000000000", -- tread, gr1
 326 => b"00011_0001_00_000101011000", -- sub, gr1, GRASS
 327 => b"00111_0000_01_000000000000", -- bne
 328 => b"00000_0000_00_000000000100", -- CONTROL_R
 329 => b"00010_1111_01_000000000000", -- add, gr15
 330 => b"00000_0000_00_000000000001", -- 1
 331 => b"00100_0000_01_000000000000", -- jump
 332 => b"00000_0000_00_000000000100", -- CONTROL_R
 333 => b"00100_0000_01_000000000000", -- jump
 334 => b"00000_0000_00_000010110011", -- COUNT_R
 335 => b"00000_0000_00_000000000000", -- 0
 336 => b"00000_0000_00_000000000000", -- 0
 337 => b"00000_0000_00_000000000000", -- 0
 338 => b"00000_0000_00_000000000000", -- 0
 339 => b"00000_0000_00_000000000000", -- 0
 340 => b"00000_0000_00_000000000000", -- 0
 341 => b"00000_0000_00_000000000000", -- 0
 342 => b"00000_0000_00_000000000000", -- 0
 343 => b"00000_0000_00_000000000001", -- 1
 344 => b"00000_0000_00_000000000000", -- 0
 345 => b"00000_0000_00_000000000001", -- 1
 346 => b"00000_0000_00_000000000010", -- 2
 347 => b"00000_0000_00_000000000011", -- 3
 348 => b"00000_0000_00_000000000100", -- 4
 349 => b"00000_0000_00_000000000000", -- 0
 350 => b"00000_0000_00_000000000000", -- 0
 351 => b"00000_0000_00_000000000000", -- 0
 352 => b"00000_0000_00_000000000000", -- 0
 353 => b"00000_0000_00_000000000000", -- 0
 354 => b"00000_0000_00_000000000000", -- 0
 355 => b"00000_0000_00_000000000000", -- 0
    



    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


