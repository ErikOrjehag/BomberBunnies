library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000010101101", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000001100011", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKBOMBS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000010", -- MAIN
  10 => b"00000_0000_00_000101001101", -- load, gr0, P1BOMBACTIVE
  11 => b"00011_0000_01_000000000000", -- sub, gr0
  12 => b"00000_0000_00_000000000001", -- 1
  13 => b"00111_0000_01_000000000000", -- bne
  14 => b"00000_0000_00_000001100001", -- TICK2
  15 => b"00000_0000_00_000101001100", -- load, gr0, P1BOMBTIME
  16 => b"00011_0000_01_000000000000", -- sub, gr0
  17 => b"00000_0000_00_000000000001", -- 1
  18 => b"00001_0000_10_000101001100", -- store, gr0, P1BOMBTIME
  19 => b"00000_0000_01_000000000000", -- load, gr0
  20 => b"00000_0000_00_000000000000", -- 0
  21 => b"00011_0000_00_000101001100", -- sub, gr0, P1BOMBTIME
  22 => b"00110_0000_01_000000000000", -- beq
  23 => b"00000_0000_00_000000011010", -- EXPLODE1
  24 => b"00100_0000_01_000000000000", -- jump
  25 => b"00000_0000_00_000001100001", -- TICK2
  26 => b"00000_0010_00_000101001011", -- load, gr2, P1BOMBPOS
  27 => b"00000_0011_00_000101010111", -- load, gr3, EXPLOSION
  28 => b"10000_0010_00_000000000000", -- tpoint, gr2
  29 => b"01110_0011_00_000000000000", -- twrite, gr3
  30 => b"00010_0010_01_000000000000", -- add, gr2
  31 => b"00000_0000_00_000000000001", -- 1
  32 => b"10000_0010_00_000000000000", -- tpoint, gr2
  33 => b"01111_0000_00_000000000000", -- tread, gr0
  34 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  35 => b"00110_0000_01_000000000000", -- beq
  36 => b"00000_0000_00_000000101110", -- P1LEFT
  37 => b"01110_0011_00_000000000000", -- twrite, gr3
  38 => b"00010_0010_01_000000000000", -- add, gr2
  39 => b"00000_0000_00_000000000001", -- 1
  40 => b"10000_0010_00_000000000000", -- tpoint, gr2
  41 => b"01111_0000_00_000000000000", -- tread, gr0
  42 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  43 => b"00110_0000_01_000000000000", -- beq
  44 => b"00000_0000_00_000000101110", -- P1LEFT
  45 => b"01110_0011_00_000000000000", -- twrite, gr3
  46 => b"00000_0010_00_000101001011", -- load, gr2, P1BOMBPOS
  47 => b"00011_0010_01_000000000000", -- sub, gr2
  48 => b"00000_0000_00_000000000001", -- 1
  49 => b"10000_0010_00_000000000000", -- tpoint, gr2
  50 => b"01111_0000_00_000000000000", -- tread, gr0
  51 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  52 => b"00110_0000_01_000000000000", -- beq
  53 => b"00000_0000_00_000000111111", -- P1DOWN
  54 => b"01110_0011_00_000000000000", -- twrite, gr3
  55 => b"00011_0010_01_000000000000", -- sub, gr2
  56 => b"00000_0000_00_000000000001", -- 1
  57 => b"10000_0010_00_000000000000", -- tpoint, gr2
  58 => b"01111_0000_00_000000000000", -- tread, gr0
  59 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  60 => b"00110_0000_01_000000000000", -- beq
  61 => b"00000_0000_00_000000111111", -- P1DOWN
  62 => b"01110_0011_00_000000000000", -- twrite, gr3
  63 => b"00000_0010_00_000101001011", -- load, gr2, P1BOMBPOS
  64 => b"00010_0010_01_000000000000", -- add, gr2
  65 => b"00000_0000_00_000000001111", -- 15
  66 => b"10000_0010_00_000000000000", -- tpoint, gr2
  67 => b"01111_0000_00_000000000000", -- tread, gr0
  68 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  69 => b"00110_0000_01_000000000000", -- beq
  70 => b"00000_0000_00_000001010000", -- P1UP
  71 => b"01110_0011_00_000000000000", -- twrite, gr3
  72 => b"00010_0010_01_000000000000", -- add, gr2
  73 => b"00000_0000_00_000000001111", -- 15
  74 => b"10000_0010_00_000000000000", -- tpoint, gr2
  75 => b"01111_0000_00_000000000000", -- tread, gr0
  76 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  77 => b"00110_0000_01_000000000000", -- beq
  78 => b"00000_0000_00_000001010000", -- P1UP
  79 => b"01110_0011_00_000000000000", -- twrite, gr3
  80 => b"00000_0010_00_000101001011", -- load, gr2, P1BOMBPOS
  81 => b"00011_0010_01_000000000000", -- sub, gr2
  82 => b"00000_0000_00_000000001111", -- 15
  83 => b"10000_0010_00_000000000000", -- tpoint, gr2
  84 => b"01111_0000_00_000000000000", -- tread, gr0
  85 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  86 => b"00110_0000_01_000000000000", -- beq
  87 => b"00000_0000_00_000001100001", -- TICK2
  88 => b"01110_0011_00_000000000000", -- twrite, gr3
  89 => b"00011_0010_01_000000000000", -- sub, gr2
  90 => b"00000_0000_00_000000001111", -- 15
  91 => b"10000_0010_00_000000000000", -- tpoint, gr2
  92 => b"01111_0000_00_000000000000", -- tread, gr0
  93 => b"00011_0000_00_000101010101", -- sub, gr0, WALL
  94 => b"00110_0000_01_000000000000", -- beq
  95 => b"00000_0000_00_000001100001", -- TICK2
  96 => b"01110_0011_00_000000000000", -- twrite, gr3
  97 => b"00100_0000_01_000000000000", -- jump
  98 => b"00000_0000_00_000000001000", -- TICKBOMBS_R
  99 => b"10101_0000_01_000000000000", -- btn1
 100 => b"00000_0000_00_000001101001", -- BTN1
 101 => b"11010_0000_01_000000000000", -- btn2
 102 => b"00000_0000_00_000010001110", -- BTN2
 103 => b"00100_0000_01_000000000000", -- jump
 104 => b"00000_0000_00_000000000110", -- BUTTON_R
 105 => b"00000_0000_00_000101010001", -- load, gr0, BOMBS1
 106 => b"00011_0000_00_000101010011", -- sub, gr0, MAXBOMBS
 107 => b"00110_0000_01_000000000000", -- beq
 108 => b"00000_0000_00_000001100101", -- BTN1_R
 109 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 110 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 111 => b"00000_0000_00_000101011010", -- load, gr0, YPOS1
 112 => b"01000_0000_01_000000000000", -- mul, gr0
 113 => b"00000_0000_00_000000001111", -- 15
 114 => b"00010_0000_00_000101011001", -- add, gr0, XPOS1
 115 => b"10000_0000_00_000000000000", -- tpoint, gr0
 116 => b"01111_0001_00_000000000000", -- tread, gr1
 117 => b"00011_0001_00_000101011000", -- sub, gr1, EGG
 118 => b"00110_0000_01_000000000000", -- beq
 119 => b"00000_0000_00_000001100111", -- BTN2_R
 120 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 121 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 122 => b"00000_0011_00_000101011010", -- load, gr3, YPOS1
 123 => b"00000_0010_00_000101011000", -- load, gr2, EGG
 124 => b"01000_0011_01_000000000000", -- mul, gr3
 125 => b"00000_0000_00_000000001111", -- 15
 126 => b"00010_0011_00_000101011001", -- add, gr3, XPOS1
 127 => b"10000_0011_00_000000000000", -- tpoint, gr3
 128 => b"01110_0010_00_000000000000", -- twrite, gr2
 129 => b"00000_0000_01_000000000000", -- load, gr0
 130 => b"00000_0000_00_000000000001", -- 1
 131 => b"00001_0000_10_000101001101", -- store, gr0, P1BOMBACTIVE
 132 => b"00001_0011_10_000101001011", -- store, gr3, P1BOMBPOS
 133 => b"00000_0000_01_000000000000", -- load, gr0
 134 => b"00000_0000_01_111101000000", -- 8000
 135 => b"00001_0000_10_000101001100", -- store, gr0, P1BOMBTIME
 136 => b"00000_0000_00_000101010001", -- load, gr0, BOMBS1
 137 => b"00010_0000_01_000000000000", -- add, gr0
 138 => b"00000_0000_00_000000000001", -- 1
 139 => b"00001_0000_10_000101010001", -- store, gr0, BOMBS1
 140 => b"00100_0000_01_000000000000", -- jump
 141 => b"00000_0000_00_000001100101", -- BTN1_R
 142 => b"00000_0000_00_000101010010", -- load, gr0, BOMBS2
 143 => b"00011_0000_00_000101010011", -- sub, gr0, MAXBOMBS
 144 => b"00110_0000_01_000000000000", -- beq
 145 => b"00000_0000_00_000001100111", -- BTN2_R
 146 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 147 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 148 => b"00000_0000_00_000101011100", -- load, gr0, YPOS2
 149 => b"01000_0000_01_000000000000", -- mul, gr0
 150 => b"00000_0000_00_000000001111", -- 15
 151 => b"00010_0000_00_000101011011", -- add, gr0, XPOS2
 152 => b"10000_0000_00_000000000000", -- tpoint, gr0
 153 => b"01111_0001_00_000000000000", -- tread, gr1
 154 => b"00011_0001_00_000101011000", -- sub, gr1, EGG
 155 => b"00110_0000_01_000000000000", -- beq
 156 => b"00000_0000_00_000001100111", -- BTN2_R
 157 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 158 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 159 => b"00000_0011_00_000101011100", -- load, gr3, YPOS2
 160 => b"00000_0010_00_000101011000", -- load, gr2, EGG
 161 => b"01000_0011_01_000000000000", -- mul, gr3
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"00010_0011_00_000101011011", -- add, gr3, XPOS2
 164 => b"10000_0011_00_000000000000", -- tpoint, gr3
 165 => b"01110_0010_00_000000000000", -- twrite, gr2
 166 => b"00000_0000_00_000101010010", -- load, gr0, BOMBS2
 167 => b"00010_0000_01_000000000000", -- add, gr0
 168 => b"00000_0000_00_000000000001", -- 1
 169 => b"00001_0000_10_000101010010", -- store, gr0, BOMBS2
 170 => b"00100_0000_01_000000000000", -- jump
 171 => b"00000_0000_00_000001100111", -- BTN2_R
 172 => b"00000_0000_00_000000000000", -- 0
 173 => b"00100_0000_01_000000000000", -- jump
 174 => b"00000_0000_00_000101001001", -- COUNT1
 175 => b"10001_0000_01_000000000000", -- joy1r
 176 => b"00000_0000_00_000011000001", -- P1R
 177 => b"10011_0000_01_000000000000", -- joy1l
 178 => b"00000_0000_00_000011100011", -- P1L
 179 => b"10010_0000_01_000000000000", -- joy1u
 180 => b"00000_0000_00_000011010010", -- P1U
 181 => b"10100_0000_01_000000000000", -- joy1d
 182 => b"00000_0000_00_000011110100", -- P1D
 183 => b"10110_0000_01_000000000000", -- joy2r
 184 => b"00000_0000_00_000100000101", -- P2R
 185 => b"11000_0000_01_000000000000", -- joy2l
 186 => b"00000_0000_00_000100100111", -- P2L
 187 => b"10111_0000_01_000000000000", -- joy2u
 188 => b"00000_0000_00_000100010110", -- P2U
 189 => b"11001_0000_01_000000000000", -- joy2d
 190 => b"00000_0000_00_000100111000", -- P2D
 191 => b"00100_0000_01_000000000000", -- jump
 192 => b"00000_0000_00_000000000100", -- CONTROL_R
 193 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 194 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 195 => b"00000_0000_00_000101011010", -- load, gr0, YPOS1
 196 => b"01000_0000_01_000000000000", -- mul, gr0
 197 => b"00000_0000_00_000000001111", -- 15
 198 => b"00010_0000_00_000101011001", -- add, gr0, XPOS1
 199 => b"00010_0000_01_000000000000", -- add, gr0
 200 => b"00000_0000_00_000000000001", -- 1
 201 => b"10000_0000_00_000000000000", -- tpoint, gr0
 202 => b"01111_0001_00_000000000000", -- tread, gr1
 203 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 204 => b"00111_0000_01_000000000000", -- bne
 205 => b"00000_0000_00_000010110011", -- J1
 206 => b"00010_1100_01_000000000000", -- add, gr12
 207 => b"00000_0000_00_000000000001", -- 1
 208 => b"00100_0000_01_000000000000", -- jump
 209 => b"00000_0000_00_000010110011", -- J1
 210 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 211 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 212 => b"00000_0000_00_000101011010", -- load, gr0, YPOS1
 213 => b"00011_0000_01_000000000000", -- sub, gr0
 214 => b"00000_0000_00_000000000001", -- 1
 215 => b"01000_0000_01_000000000000", -- mul, gr0
 216 => b"00000_0000_00_000000001111", -- 15
 217 => b"00010_0000_00_000101011001", -- add, gr0, XPOS1
 218 => b"10000_0000_00_000000000000", -- tpoint, gr0
 219 => b"01111_0001_00_000000000000", -- tread, gr1
 220 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 221 => b"00111_0000_01_000000000000", -- bne
 222 => b"00000_0000_00_000010110111", -- J2
 223 => b"00011_1101_01_000000000000", -- sub, gr13
 224 => b"00000_0000_00_000000000001", -- 1
 225 => b"00100_0000_01_000000000000", -- jump
 226 => b"00000_0000_00_000010110111", -- J2
 227 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 228 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 229 => b"00000_0000_00_000101011010", -- load, gr0, YPOS1
 230 => b"01000_0000_01_000000000000", -- mul, gr0
 231 => b"00000_0000_00_000000001111", -- 15
 232 => b"00010_0000_00_000101011001", -- add, gr0, XPOS1
 233 => b"00011_0000_01_000000000000", -- sub, gr0
 234 => b"00000_0000_00_000000000001", -- 1
 235 => b"10000_0000_00_000000000000", -- tpoint, gr0
 236 => b"01111_0001_00_000000000000", -- tread, gr1
 237 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 238 => b"00111_0000_01_000000000000", -- bne
 239 => b"00000_0000_00_000010110011", -- J1
 240 => b"00011_1100_01_000000000000", -- sub, gr12
 241 => b"00000_0000_00_000000000001", -- 1
 242 => b"00100_0000_01_000000000000", -- jump
 243 => b"00000_0000_00_000010110011", -- J1
 244 => b"00001_1100_10_000101011001", -- store, gr12, XPOS1
 245 => b"00001_1101_10_000101011010", -- store, gr13, YPOS1
 246 => b"00000_0000_00_000101011010", -- load, gr0, YPOS1
 247 => b"00010_0000_01_000000000000", -- add, gr0
 248 => b"00000_0000_00_000000000001", -- 1
 249 => b"01000_0000_01_000000000000", -- mul, gr0
 250 => b"00000_0000_00_000000001111", -- 15
 251 => b"00010_0000_00_000101011001", -- add, gr0, XPOS1
 252 => b"10000_0000_00_000000000000", -- tpoint, gr0
 253 => b"01111_0001_00_000000000000", -- tread, gr1
 254 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 255 => b"00111_0000_01_000000000000", -- bne
 256 => b"00000_0000_00_000010110111", -- J2
 257 => b"00010_1101_01_000000000000", -- add, gr13
 258 => b"00000_0000_00_000000000001", -- 1
 259 => b"00100_0000_01_000000000000", -- jump
 260 => b"00000_0000_00_000010110111", -- J2
 261 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 262 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 263 => b"00000_0000_00_000101011100", -- load, gr0, YPOS2
 264 => b"01000_0000_01_000000000000", -- mul, gr0
 265 => b"00000_0000_00_000000001111", -- 15
 266 => b"00010_0000_00_000101011011", -- add, gr0, XPOS2
 267 => b"00010_0000_01_000000000000", -- add, gr0
 268 => b"00000_0000_00_000000000001", -- 1
 269 => b"10000_0000_00_000000000000", -- tpoint, gr0
 270 => b"01111_0001_00_000000000000", -- tread, gr1
 271 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 272 => b"00111_0000_01_000000000000", -- bne
 273 => b"00000_0000_00_000010111011", -- J3
 274 => b"00010_1110_01_000000000000", -- add, gr14
 275 => b"00000_0000_00_000000000001", -- 1
 276 => b"00100_0000_01_000000000000", -- jump
 277 => b"00000_0000_00_000010111011", -- J3
 278 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 279 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 280 => b"00000_0000_00_000101011100", -- load, gr0, YPOS2
 281 => b"00011_0000_01_000000000000", -- sub, gr0
 282 => b"00000_0000_00_000000000001", -- 1
 283 => b"01000_0000_01_000000000000", -- mul, gr0
 284 => b"00000_0000_00_000000001111", -- 15
 285 => b"00010_0000_00_000101011011", -- add, gr0, XPOS2
 286 => b"10000_0000_00_000000000000", -- tpoint, gr0
 287 => b"01111_0001_00_000000000000", -- tread, gr1
 288 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 289 => b"00111_0000_01_000000000000", -- bne
 290 => b"00000_0000_00_000000000100", -- CONTROL_R
 291 => b"00011_1111_01_000000000000", -- sub, gr15
 292 => b"00000_0000_00_000000000001", -- 1
 293 => b"00100_0000_01_000000000000", -- jump
 294 => b"00000_0000_00_000000000100", -- CONTROL_R
 295 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 296 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 297 => b"00000_0000_00_000101011100", -- load, gr0, YPOS2
 298 => b"01000_0000_01_000000000000", -- mul, gr0
 299 => b"00000_0000_00_000000001111", -- 15
 300 => b"00010_0000_00_000101011011", -- add, gr0, XPOS2
 301 => b"00011_0000_01_000000000000", -- sub, gr0
 302 => b"00000_0000_00_000000000001", -- 1
 303 => b"10000_0000_00_000000000000", -- tpoint, gr0
 304 => b"01111_0001_00_000000000000", -- tread, gr1
 305 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 306 => b"00111_0000_01_000000000000", -- bne
 307 => b"00000_0000_00_000010111011", -- J3
 308 => b"00011_1110_01_000000000000", -- sub, gr14
 309 => b"00000_0000_00_000000000001", -- 1
 310 => b"00100_0000_01_000000000000", -- jump
 311 => b"00000_0000_00_000010111011", -- J3
 312 => b"00001_1110_10_000101011011", -- store, gr14, XPOS2
 313 => b"00001_1111_10_000101011100", -- store, gr15, YPOS2
 314 => b"00000_0000_00_000101011100", -- load, gr0, YPOS2
 315 => b"00010_0000_01_000000000000", -- add, gr0
 316 => b"00000_0000_00_000000000001", -- 1
 317 => b"01000_0000_01_000000000000", -- mul, gr0
 318 => b"00000_0000_00_000000001111", -- 15
 319 => b"00010_0000_00_000101011011", -- add, gr0, XPOS2
 320 => b"10000_0000_00_000000000000", -- tpoint, gr0
 321 => b"01111_0001_00_000000000000", -- tread, gr1
 322 => b"00011_0001_00_000101010100", -- sub, gr1, GRASS
 323 => b"00111_0000_01_000000000000", -- bne
 324 => b"00000_0000_00_000000000100", -- CONTROL_R
 325 => b"00010_1111_01_000000000000", -- add, gr15
 326 => b"00000_0000_00_000000000001", -- 1
 327 => b"00100_0000_01_000000000000", -- jump
 328 => b"00000_0000_00_000000000100", -- CONTROL_R
 329 => b"00100_0000_01_000000000000", -- jump
 330 => b"00000_0000_00_000010101111", -- COUNT_R
 331 => b"00000_0000_00_000000000000", -- 0
 332 => b"00000_0000_00_000000000000", -- 0
 333 => b"00000_0000_00_000000000000", -- 0
 334 => b"00000_0000_00_000000000000", -- 0
 335 => b"00000_0000_00_000000000000", -- 0
 336 => b"00000_0000_00_000000000000", -- 0
 337 => b"00000_0000_00_000000000000", -- 0
 338 => b"00000_0000_00_000000000000", -- 0
 339 => b"00000_0000_00_000000000001", -- 1
 340 => b"00000_0000_00_000000000000", -- 0
 341 => b"00000_0000_00_000000000001", -- 1
 342 => b"00000_0000_00_000000000010", -- 2
 343 => b"00000_0000_00_000000000011", -- 3
 344 => b"00000_0000_00_000000000100", -- 4
 345 => b"00000_0000_00_000000000000", -- 0
 346 => b"00000_0000_00_000000000000", -- 0
 347 => b"00000_0000_00_000000000000", -- 0
 348 => b"00000_0000_00_000000000000", -- 0
 349 => b"00000_0000_00_000000000000", -- 0
 350 => b"00000_0000_00_000000000000", -- 0
 351 => b"00000_0000_00_000000000000", -- 0


    others => (others => 0)
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = 1 then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = 1 else PM(to_integer(pAddr));

end Behavioral; 
