library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_0000_01_000000000000", -- load, gr0
   1 => b"00000_0000_00_000000000000", -- 0
   2 => b"00001_0000_10_010001011100", -- store, gr0, P1DEAD
   3 => b"00001_0000_10_010001011101", -- store, gr0, P2DEAD
   4 => b"00001_0000_10_010010000100", -- store, gr0, P1BOMBCOUNT
   5 => b"00001_0000_10_010010000101", -- store, gr0, P2BOMBCOUNT
   6 => b"00000_1100_01_000000000000", -- load, gr12
   7 => b"00000_0000_00_000000000001", -- 1
   8 => b"00000_1101_01_000000000000", -- load, gr13
   9 => b"00000_0000_00_000000000001", -- 1
  10 => b"00000_1110_01_000000000000", -- load, gr14
  11 => b"00000_0000_00_000000001101", -- 13
  12 => b"00000_1111_01_000000000000", -- load, gr15
  13 => b"00000_0000_00_000000001011", -- 11
  14 => b"00001_0000_10_010001100000", -- store, gr0, P1BOMB1POS
  15 => b"00001_0000_10_010001100010", -- store, gr0, P1BOMB1ACTIVE
  16 => b"00001_0000_10_010001100001", -- store, gr0, P1BOMB1TIME
  17 => b"00001_0000_10_010001100110", -- store, gr0, P1BOMB2POS
  18 => b"00001_0000_10_010001101000", -- store, gr0, P1BOMB2ACTIVE
  19 => b"00001_0000_10_010001100111", -- store, gr0, P1BOMB2TIME
  20 => b"00001_0000_10_010001101100", -- store, gr0, P1BOMB3POS
  21 => b"00001_0000_10_010001101110", -- store, gr0, P1BOMB3ACTIVE
  22 => b"00001_0000_10_010001101101", -- store, gr0, P1BOMB3TIME
  23 => b"00001_0000_10_010001110010", -- store, gr0, P2BOMB1POS
  24 => b"00001_0000_10_010001110100", -- store, gr0, P2BOMB1ACTIVE
  25 => b"00001_0000_10_010001110011", -- store, gr0, P2BOMB1TIME
  26 => b"00001_0000_10_010001111000", -- store, gr0, P2BOMB2POS
  27 => b"00001_0000_10_010001111010", -- store, gr0, P2BOMB2ACTIVE
  28 => b"00001_0000_10_010001111001", -- store, gr0, P2BOMB2TIME
  29 => b"00001_0000_10_010001111110", -- store, gr0, P2BOMB3POS
  30 => b"00001_0000_10_010010000000", -- store, gr0, P2BOMB3ACTIVE
  31 => b"00001_0000_10_010001111111", -- store, gr0, P2BOMB3TIME
  32 => b"00001_0000_10_010001100101", -- store, gr0, P1EXPLOSION1POS
  33 => b"00001_0000_10_010001100100", -- store, gr0, P1EXPLOSION1ACTIVE
  34 => b"00001_0000_10_010001100011", -- store, gr0, P1EXPLOSION1TIME
  35 => b"00001_0000_10_010001101011", -- store, gr0, P1EXPLOSION2POS
  36 => b"00001_0000_10_010001101010", -- store, gr0, P1EXPLOSION2ACTIVE
  37 => b"00001_0000_10_010001101001", -- store, gr0, P1EXPLOSION2TIME
  38 => b"00001_0000_10_010001110001", -- store, gr0, P1EXPLOSION3POS
  39 => b"00001_0000_10_010001110000", -- store, gr0, P1EXPLOSION3ACTIVE
  40 => b"00001_0000_10_010001101111", -- store, gr0, P1EXPLOSION3TIME
  41 => b"00001_0000_10_010001110111", -- store, gr0, P2EXPLOSION1POS
  42 => b"00001_0000_10_010001110110", -- store, gr0, P2EXPLOSION1ACTIVE
  43 => b"00001_0000_10_010001110101", -- store, gr0, P2EXPLOSION1TIME
  44 => b"00001_0000_10_010001111101", -- store, gr0, P2EXPLOSION2POS
  45 => b"00001_0000_10_010001111100", -- store, gr0, P2EXPLOSION2ACTIVE
  46 => b"00001_0000_10_010001111011", -- store, gr0, P2EXPLOSION2TIME
  47 => b"00001_0000_10_010010000011", -- store, gr0, P2EXPLOSION3POS
  48 => b"00001_0000_10_010010000010", -- store, gr0, P2EXPLOSION3ACTIVE
  49 => b"00001_0000_10_010010000001", -- store, gr0, P2EXPLOSION3TIME
  50 => b"00000_0000_01_000000000000", -- load, gr0
  51 => b"00000_0000_00_000000000000", -- 0
  52 => b"00000_0011_01_000000000000", -- load, gr3
  53 => b"00000_0000_00_000011000011", -- 195
  54 => b"00001_0000_10_010010001011", -- store, gr0, MOVE
  55 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
  56 => b"00001_0011_10_010010001011", -- store, gr3, MOVE
  57 => b"00011_0010_00_010010001011", -- sub, gr2, MOVE
  58 => b"00110_0000_01_000000000000", -- beq
  59 => b"00000_0000_00_000001000111", -- INITEND
  60 => b"10000_0000_00_000000000000", -- tpoint, gr0
  61 => b"01111_0001_00_000000000000", -- tread, gr1
  62 => b"00011_0001_00_010010001111", -- sub, gr1, WALL
  63 => b"00110_0000_01_000000000000", -- beq
  64 => b"00000_0000_00_000001000011", -- INCREASE
  65 => b"00000_0001_00_010010010000", -- load, gr1, BREAKABLE
  66 => b"01110_0001_00_000000000000", -- twrite, gr1
  67 => b"00010_0000_01_000000000000", -- add, gr0
  68 => b"00000_0000_00_000000000001", -- 1
  69 => b"00100_0000_01_000000000000", -- jump
  70 => b"00000_0000_00_000000110110", -- INITLOOP
  71 => b"00000_0000_00_010010001110", -- load, gr0, GRASS
  72 => b"00000_0001_01_000000000000", -- load, gr1
  73 => b"00000_0000_00_000000010000", -- 16
  74 => b"10000_0001_00_000000000000", -- tpoint, gr1
  75 => b"01110_0000_00_000000000000", -- twrite, gr0
  76 => b"00010_0001_01_000000000000", -- add, gr1
  77 => b"00000_0000_00_000000000001", -- 1
  78 => b"10000_0001_00_000000000000", -- tpoint, gr1
  79 => b"01110_0000_00_000000000000", -- twrite, gr0
  80 => b"00010_0001_01_000000000000", -- add, gr1
  81 => b"00000_0000_00_000000001110", -- 14
  82 => b"10000_0001_00_000000000000", -- tpoint, gr1
  83 => b"01110_0000_00_000000000000", -- twrite, gr0
  84 => b"00000_0001_01_000000000000", -- load, gr1
  85 => b"00000_0000_00_000010110010", -- 178
  86 => b"10000_0001_00_000000000000", -- tpoint, gr1
  87 => b"01110_0000_00_000000000000", -- twrite, gr0
  88 => b"00011_0001_01_000000000000", -- sub, gr1
  89 => b"00000_0000_00_000000000001", -- 1
  90 => b"10000_0001_00_000000000000", -- tpoint, gr1
  91 => b"01110_0000_00_000000000000", -- twrite, gr0
  92 => b"00011_0001_01_000000000000", -- sub, gr1
  93 => b"00000_0000_00_000000001110", -- 14
  94 => b"10000_0001_00_000000000000", -- tpoint, gr1
  95 => b"01110_0000_00_000000000000", -- twrite, gr0
  96 => b"00100_0000_01_000000000000", -- jump
  97 => b"00000_0000_00_000010101000", -- CHECKDEATH
  98 => b"00100_0000_01_000000000000", -- jump
  99 => b"00000_0000_00_000001101110", -- CHECKBOMBDEATH
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_001110111000", -- CONTROL
 102 => b"00100_0000_01_000000000000", -- jump
 103 => b"00000_0000_00_001011110010", -- BUTTON
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000111001111", -- TICKBOMBS
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 108 => b"00100_0000_01_000000000000", -- jump
 109 => b"00000_0000_00_000001100000", -- MAIN
 110 => b"00000_0010_01_000000000000", -- load, gr2
 111 => b"00000_0000_00_000000000001", -- 1
 112 => b"00000_0000_00_010001100000", -- load, gr0, P1BOMB1POS
 113 => b"10000_0000_00_000000000000", -- tpoint, gr0
 114 => b"01111_0001_00_000000000000", -- tread, gr1
 115 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 116 => b"00110_0000_01_000000000000", -- beq
 117 => b"00000_0000_00_000010010110", -- P1BOMB1DETONATE
 118 => b"00000_0000_00_010001100110", -- load, gr0, P1BOMB2POS
 119 => b"10000_0000_00_000000000000", -- tpoint, gr0
 120 => b"01111_0001_00_000000000000", -- tread, gr1
 121 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 122 => b"00110_0000_01_000000000000", -- beq
 123 => b"00000_0000_00_000010011001", -- P1BOMB2DETONATE
 124 => b"00000_0000_00_010001101100", -- load, gr0, P1BOMB3POS
 125 => b"10000_0000_00_000000000000", -- tpoint, gr0
 126 => b"01111_0001_00_000000000000", -- tread, gr1
 127 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 128 => b"00110_0000_01_000000000000", -- beq
 129 => b"00000_0000_00_000010011100", -- P1BOMB3DETONATE
 130 => b"00000_0000_00_010001110010", -- load, gr0, P2BOMB1POS
 131 => b"10000_0000_00_000000000000", -- tpoint, gr0
 132 => b"01111_0001_00_000000000000", -- tread, gr1
 133 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 134 => b"00110_0000_01_000000000000", -- beq
 135 => b"00000_0000_00_000010011111", -- P2BOMB1DETONATE
 136 => b"00000_0000_00_010001111000", -- load, gr0, P2BOMB2POS
 137 => b"10000_0000_00_000000000000", -- tpoint, gr0
 138 => b"01111_0001_00_000000000000", -- tread, gr1
 139 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 140 => b"00110_0000_01_000000000000", -- beq
 141 => b"00000_0000_00_000010100010", -- P2BOMB2DETONATE
 142 => b"00000_0000_00_010001111110", -- load, gr0, P2BOMB3POS
 143 => b"10000_0000_00_000000000000", -- tpoint, gr0
 144 => b"01111_0001_00_000000000000", -- tread, gr1
 145 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 146 => b"00110_0000_01_000000000000", -- beq
 147 => b"00000_0000_00_000010100101", -- P2BOMB3DETONATE
 148 => b"00100_0000_01_000000000000", -- jump
 149 => b"00000_0000_00_000001100100", -- CHECKBOMBDEATH_R
 150 => b"00001_0010_10_010001100001", -- store, gr2, P1BOMB1TIME
 151 => b"00100_0000_01_000000000000", -- jump
 152 => b"00000_0000_00_000001110110", -- P1BOMB1DETONATE_R
 153 => b"00001_0010_10_010001100111", -- store, gr2, P1BOMB2TIME
 154 => b"00100_0000_01_000000000000", -- jump
 155 => b"00000_0000_00_000001111100", -- P1BOMB2DETONATE_R
 156 => b"00001_0010_10_010001101101", -- store, gr2, P1BOMB3TIME
 157 => b"00100_0000_01_000000000000", -- jump
 158 => b"00000_0000_00_000010000010", -- P1BOMB3DETONATE_R
 159 => b"00001_0010_10_010001110011", -- store, gr2, P2BOMB1TIME
 160 => b"00100_0000_01_000000000000", -- jump
 161 => b"00000_0000_00_000010001000", -- P2BOMB1DETONATE_R
 162 => b"00001_0010_10_010001111001", -- store, gr2, P2BOMB2TIME
 163 => b"00100_0000_01_000000000000", -- jump
 164 => b"00000_0000_00_000010001110", -- P2BOMB2DETONATE_R
 165 => b"00001_0010_10_010001111111", -- store, gr2, P2BOMB3TIME
 166 => b"00100_0000_01_000000000000", -- jump
 167 => b"00000_0000_00_000010010100", -- P2BOMB3DETONATE_R
 168 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 169 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 170 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 171 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 172 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
 173 => b"01000_0000_01_000000000000", -- mul, gr0
 174 => b"00000_0000_00_000000001111", -- 15
 175 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
 176 => b"10000_0000_00_000000000000", -- tpoint, gr0
 177 => b"01111_0001_00_000000000000", -- tread, gr1
 178 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 179 => b"00110_0000_01_000000000000", -- beq
 180 => b"00000_0000_00_000011000000", -- P1DEATH
 181 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
 182 => b"01000_0000_01_000000000000", -- mul, gr0
 183 => b"00000_0000_00_000000001111", -- 15
 184 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
 185 => b"10000_0000_00_000000000000", -- tpoint, gr0
 186 => b"01111_0001_00_000000000000", -- tread, gr1
 187 => b"00011_0001_00_010010010001", -- sub, gr1, EXPLOSION
 188 => b"00110_0000_01_000000000000", -- beq
 189 => b"00000_0000_00_000011010100", -- P2DEATH
 190 => b"00100_0000_01_000000000000", -- jump
 191 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 192 => b"00000_0000_01_000000000000", -- load, gr0
 193 => b"00000_0000_00_000000000001", -- 1
 194 => b"00001_0000_10_010001011100", -- store, gr0, P1DEAD
 195 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 196 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 197 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
 198 => b"01000_0000_01_000000000000", -- mul, gr0
 199 => b"00000_0000_00_000000001111", -- 15
 200 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
 201 => b"00001_0000_10_010001011110", -- store, gr0, DEADPOS1
 202 => b"10000_0000_00_000000000000", -- tpoint, gr0
 203 => b"00000_0000_01_000000000000", -- load, gr0
 204 => b"00000_0000_00_000000000101", -- 5
 205 => b"01110_0000_00_000000000000", -- twrite, gr0
 206 => b"00000_1100_01_000000000000", -- load, gr12
 207 => b"00000_0000_00_000000000000", -- 0
 208 => b"00000_1101_01_000000000000", -- load, gr13
 209 => b"00000_0000_00_000000010000", -- 16
 210 => b"00100_0000_01_000000000000", -- jump
 211 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 212 => b"00000_0000_01_000000000000", -- load, gr0
 213 => b"00000_0000_00_000000000001", -- 1
 214 => b"00001_0000_10_010001011101", -- store, gr0, P2DEAD
 215 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 216 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 217 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
 218 => b"01000_0000_01_000000000000", -- mul, gr0
 219 => b"00000_0000_00_000000001111", -- 15
 220 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
 221 => b"00001_0000_10_010001011111", -- store, gr0, DEADPOS2
 222 => b"10000_0000_00_000000000000", -- tpoint, gr0
 223 => b"00000_0000_01_000000000000", -- load, gr0
 224 => b"00000_0000_00_000000000101", -- 5
 225 => b"01110_0000_00_000000000000", -- twrite, gr0
 226 => b"00000_1110_01_000000000000", -- load, gr14
 227 => b"00000_0000_00_000000000000", -- 0
 228 => b"00000_1111_01_000000000000", -- load, gr15
 229 => b"00000_0000_00_000000010000", -- 16
 230 => b"00100_0000_01_000000000000", -- jump
 231 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 232 => b"00000_0000_00_010001100100", -- load, gr0, P1EXPLOSION1ACTIVE
 233 => b"00011_0000_01_000000000000", -- sub, gr0
 234 => b"00000_0000_00_000000000001", -- 1
 235 => b"00111_0000_01_000000000000", -- bne
 236 => b"00000_0000_00_000011110110", -- P1EXPLOSION2
 237 => b"00000_0000_00_010001100011", -- load, gr0, P1EXPLOSION1TIME
 238 => b"00011_0000_01_000000000000", -- sub, gr0
 239 => b"00000_0000_00_000000000001", -- 1
 240 => b"00001_0000_10_010001100011", -- store, gr0, P1EXPLOSION1TIME
 241 => b"00000_0000_01_000000000000", -- load, gr0
 242 => b"00000_0000_00_000000000000", -- 0
 243 => b"00011_0000_00_010001100011", -- sub, gr0, P1EXPLOSION1TIME
 244 => b"00110_0000_01_000000000000", -- beq
 245 => b"00000_0000_00_000100111110", -- P1EXPLOSION1FADE
 246 => b"00000_0000_00_010001101010", -- load, gr0, P1EXPLOSION2ACTIVE
 247 => b"00011_0000_01_000000000000", -- sub, gr0
 248 => b"00000_0000_00_000000000001", -- 1
 249 => b"00111_0000_01_000000000000", -- bne
 250 => b"00000_0000_00_000100000100", -- P1EXPLOSION3
 251 => b"00000_0000_00_010001101001", -- load, gr0, P1EXPLOSION2TIME
 252 => b"00011_0000_01_000000000000", -- sub, gr0
 253 => b"00000_0000_00_000000000001", -- 1
 254 => b"00001_0000_10_010001101001", -- store, gr0, P1EXPLOSION2TIME
 255 => b"00000_0000_01_000000000000", -- load, gr0
 256 => b"00000_0000_00_000000000000", -- 0
 257 => b"00011_0000_00_010001101001", -- sub, gr0, P1EXPLOSION2TIME
 258 => b"00110_0000_01_000000000000", -- beq
 259 => b"00000_0000_00_000101000100", -- P1EXPLOSION2FADE
 260 => b"00000_0000_00_010001110000", -- load, gr0, P1EXPLOSION3ACTIVE
 261 => b"00011_0000_01_000000000000", -- sub, gr0
 262 => b"00000_0000_00_000000000001", -- 1
 263 => b"00111_0000_01_000000000000", -- bne
 264 => b"00000_0000_00_000100010010", -- P2EXPLOSION1
 265 => b"00000_0000_00_010001101111", -- load, gr0, P1EXPLOSION3TIME
 266 => b"00011_0000_01_000000000000", -- sub, gr0
 267 => b"00000_0000_00_000000000001", -- 1
 268 => b"00001_0000_10_010001101111", -- store, gr0, P1EXPLOSION3TIME
 269 => b"00000_0000_01_000000000000", -- load, gr0
 270 => b"00000_0000_00_000000000000", -- 0
 271 => b"00011_0000_00_010001101111", -- sub, gr0, P1EXPLOSION3TIME
 272 => b"00110_0000_01_000000000000", -- beq
 273 => b"00000_0000_00_000101001010", -- P1EXPLOSION3FADE
 274 => b"00000_0000_00_010001110110", -- load, gr0, P2EXPLOSION1ACTIVE
 275 => b"00011_0000_01_000000000000", -- sub, gr0
 276 => b"00000_0000_00_000000000001", -- 1
 277 => b"00111_0000_01_000000000000", -- bne
 278 => b"00000_0000_00_000100100000", -- P2EXPLOSION2
 279 => b"00000_0000_00_010001110101", -- load, gr0, P2EXPLOSION1TIME
 280 => b"00011_0000_01_000000000000", -- sub, gr0
 281 => b"00000_0000_00_000000000001", -- 1
 282 => b"00001_0000_10_010001110101", -- store, gr0, P2EXPLOSION1TIME
 283 => b"00000_0000_01_000000000000", -- load, gr0
 284 => b"00000_0000_00_000000000000", -- 0
 285 => b"00011_0000_00_010001110101", -- sub, gr0, P2EXPLOSION1TIME
 286 => b"00110_0000_01_000000000000", -- beq
 287 => b"00000_0000_00_000101010000", -- P2EXPLOSION1FADE
 288 => b"00000_0000_00_010001111100", -- load, gr0, P2EXPLOSION2ACTIVE
 289 => b"00011_0000_01_000000000000", -- sub, gr0
 290 => b"00000_0000_00_000000000001", -- 1
 291 => b"00111_0000_01_000000000000", -- bne
 292 => b"00000_0000_00_000100101110", -- P2EXPLOSION3
 293 => b"00000_0000_00_010001111011", -- load, gr0, P2EXPLOSION2TIME
 294 => b"00011_0000_01_000000000000", -- sub, gr0
 295 => b"00000_0000_00_000000000001", -- 1
 296 => b"00001_0000_10_010001111011", -- store, gr0, P2EXPLOSION2TIME
 297 => b"00000_0000_01_000000000000", -- load, gr0
 298 => b"00000_0000_00_000000000000", -- 0
 299 => b"00011_0000_00_010001111011", -- sub, gr0, P2EXPLOSION2TIME
 300 => b"00110_0000_01_000000000000", -- beq
 301 => b"00000_0000_00_000101010110", -- P2EXPLOSION2FADE
 302 => b"00000_0000_00_010010000010", -- load, gr0, P2EXPLOSION3ACTIVE
 303 => b"00011_0000_01_000000000000", -- sub, gr0
 304 => b"00000_0000_00_000000000001", -- 1
 305 => b"00111_0000_01_000000000000", -- bne
 306 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 307 => b"00000_0000_00_010010000001", -- load, gr0, P2EXPLOSION3TIME
 308 => b"00011_0000_01_000000000000", -- sub, gr0
 309 => b"00000_0000_00_000000000001", -- 1
 310 => b"00001_0000_10_010010000001", -- store, gr0, P2EXPLOSION3TIME
 311 => b"00000_0000_01_000000000000", -- load, gr0
 312 => b"00000_0000_00_000000000000", -- 0
 313 => b"00011_0000_00_010010000001", -- sub, gr0, P2EXPLOSION3TIME
 314 => b"00110_0000_01_000000000000", -- beq
 315 => b"00000_0000_00_000101011100", -- P2EXPLOSION3FADE
 316 => b"00100_0000_01_000000000000", -- jump
 317 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 318 => b"00000_0000_01_000000000000", -- load, gr0
 319 => b"00000_0000_00_000000000000", -- 0
 320 => b"00001_0000_10_010001100100", -- store, gr0, P1EXPLOSION1ACTIVE
 321 => b"00000_0100_00_010001100101", -- load, gr4, P1EXPLOSION1POS
 322 => b"00100_0000_01_000000000000", -- jump
 323 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 324 => b"00000_0000_01_000000000000", -- load, gr0
 325 => b"00000_0000_00_000000000000", -- 0
 326 => b"00001_0000_10_010001101010", -- store, gr0, P1EXPLOSION2ACTIVE
 327 => b"00000_0100_00_010001101011", -- load, gr4, P1EXPLOSION2POS
 328 => b"00100_0000_01_000000000000", -- jump
 329 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 330 => b"00000_0000_01_000000000000", -- load, gr0
 331 => b"00000_0000_00_000000000000", -- 0
 332 => b"00001_0000_10_010001110000", -- store, gr0, P1EXPLOSION3ACTIVE
 333 => b"00000_0100_00_010001110001", -- load, gr4, P1EXPLOSION3POS
 334 => b"00100_0000_01_000000000000", -- jump
 335 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 336 => b"00000_0000_01_000000000000", -- load, gr0
 337 => b"00000_0000_00_000000000000", -- 0
 338 => b"00001_0000_10_010001110110", -- store, gr0, P2EXPLOSION1ACTIVE
 339 => b"00000_0100_00_010001110111", -- load, gr4, P2EXPLOSION1POS
 340 => b"00100_0000_01_000000000000", -- jump
 341 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 342 => b"00000_0000_01_000000000000", -- load, gr0
 343 => b"00000_0000_00_000000000000", -- 0
 344 => b"00001_0000_10_010001111100", -- store, gr0, P2EXPLOSION2ACTIVE
 345 => b"00000_0100_00_010001111101", -- load, gr4, P2EXPLOSION2POS
 346 => b"00100_0000_01_000000000000", -- jump
 347 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 348 => b"00000_0000_01_000000000000", -- load, gr0
 349 => b"00000_0000_00_000000000000", -- 0
 350 => b"00001_0000_10_010010000010", -- store, gr0, P2EXPLOSION3ACTIVE
 351 => b"00000_0100_00_010010000011", -- load, gr4, P2EXPLOSION3POS
 352 => b"00100_0000_01_000000000000", -- jump
 353 => b"00000_0000_00_000101100010", -- FADEEXPLOSION
 354 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 355 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 356 => b"00000_0011_00_010010001110", -- load, gr3, GRASS
 357 => b"10000_0010_00_000000000000", -- tpoint, gr2
 358 => b"01110_0011_00_000000000000", -- twrite, gr3
 359 => b"00010_0010_01_000000000000", -- add, gr2
 360 => b"00000_0000_00_000000000001", -- 1
 361 => b"10000_0010_00_000000000000", -- tpoint, gr2
 362 => b"01111_0000_00_000000000000", -- tread, gr0
 363 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 364 => b"00110_0000_01_000000000000", -- beq
 365 => b"00000_0000_00_000101111111", -- FADELEFT
 366 => b"01111_0000_00_000000000000", -- tread, gr0
 367 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 368 => b"00110_0000_01_000000000000", -- beq
 369 => b"00000_0000_00_000101111111", -- FADELEFT
 370 => b"01110_0011_00_000000000000", -- twrite, gr3
 371 => b"00010_0010_01_000000000000", -- add, gr2
 372 => b"00000_0000_00_000000000001", -- 1
 373 => b"10000_0010_00_000000000000", -- tpoint, gr2
 374 => b"01111_0000_00_000000000000", -- tread, gr0
 375 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 376 => b"00110_0000_01_000000000000", -- beq
 377 => b"00000_0000_00_000101111111", -- FADELEFT
 378 => b"01111_0000_00_000000000000", -- tread, gr0
 379 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 380 => b"00110_0000_01_000000000000", -- beq
 381 => b"00000_0000_00_000101111111", -- FADELEFT
 382 => b"01110_0011_00_000000000000", -- twrite, gr3
 383 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 384 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 385 => b"00011_0010_01_000000000000", -- sub, gr2
 386 => b"00000_0000_00_000000000001", -- 1
 387 => b"10000_0010_00_000000000000", -- tpoint, gr2
 388 => b"01111_0000_00_000000000000", -- tread, gr0
 389 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 390 => b"00110_0000_01_000000000000", -- beq
 391 => b"00000_0000_00_000110011001", -- FADEDOWN
 392 => b"01111_0000_00_000000000000", -- tread, gr0
 393 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 394 => b"00110_0000_01_000000000000", -- beq
 395 => b"00000_0000_00_000110011001", -- FADEDOWN
 396 => b"01110_0011_00_000000000000", -- twrite, gr3
 397 => b"00011_0010_01_000000000000", -- sub, gr2
 398 => b"00000_0000_00_000000000001", -- 1
 399 => b"10000_0010_00_000000000000", -- tpoint, gr2
 400 => b"01111_0000_00_000000000000", -- tread, gr0
 401 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 402 => b"00110_0000_01_000000000000", -- beq
 403 => b"00000_0000_00_000110011001", -- FADEDOWN
 404 => b"01111_0000_00_000000000000", -- tread, gr0
 405 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 406 => b"00110_0000_01_000000000000", -- beq
 407 => b"00000_0000_00_000110011001", -- FADEDOWN
 408 => b"01110_0011_00_000000000000", -- twrite, gr3
 409 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 410 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 411 => b"00010_0010_01_000000000000", -- add, gr2
 412 => b"00000_0000_00_000000001111", -- 15
 413 => b"10000_0010_00_000000000000", -- tpoint, gr2
 414 => b"01111_0000_00_000000000000", -- tread, gr0
 415 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 416 => b"00110_0000_01_000000000000", -- beq
 417 => b"00000_0000_00_000110110011", -- FADEUP
 418 => b"01111_0000_00_000000000000", -- tread, gr0
 419 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 420 => b"00110_0000_01_000000000000", -- beq
 421 => b"00000_0000_00_000110110011", -- FADEUP
 422 => b"01110_0011_00_000000000000", -- twrite, gr3
 423 => b"00010_0010_01_000000000000", -- add, gr2
 424 => b"00000_0000_00_000000001111", -- 15
 425 => b"10000_0010_00_000000000000", -- tpoint, gr2
 426 => b"01111_0000_00_000000000000", -- tread, gr0
 427 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 428 => b"00110_0000_01_000000000000", -- beq
 429 => b"00000_0000_00_000110110011", -- FADEUP
 430 => b"01111_0000_00_000000000000", -- tread, gr0
 431 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 432 => b"00110_0000_01_000000000000", -- beq
 433 => b"00000_0000_00_000110110011", -- FADEUP
 434 => b"01110_0011_00_000000000000", -- twrite, gr3
 435 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 436 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 437 => b"00011_0010_01_000000000000", -- sub, gr2
 438 => b"00000_0000_00_000000001111", -- 15
 439 => b"10000_0010_00_000000000000", -- tpoint, gr2
 440 => b"01111_0000_00_000000000000", -- tread, gr0
 441 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 442 => b"00110_0000_01_000000000000", -- beq
 443 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 444 => b"01111_0000_00_000000000000", -- tread, gr0
 445 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 446 => b"00110_0000_01_000000000000", -- beq
 447 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 448 => b"01110_0011_00_000000000000", -- twrite, gr3
 449 => b"00011_0010_01_000000000000", -- sub, gr2
 450 => b"00000_0000_00_000000001111", -- 15
 451 => b"10000_0010_00_000000000000", -- tpoint, gr2
 452 => b"01111_0000_00_000000000000", -- tread, gr0
 453 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 454 => b"00110_0000_01_000000000000", -- beq
 455 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 456 => b"01111_0000_00_000000000000", -- tread, gr0
 457 => b"00011_0000_00_010010010000", -- sub, gr0, BREAKABLE
 458 => b"00110_0000_01_000000000000", -- beq
 459 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 460 => b"01110_0011_00_000000000000", -- twrite, gr3
 461 => b"00100_0000_01_000000000000", -- jump
 462 => b"00000_0000_00_000011101000", -- TICKEXPLOSIONS
 463 => b"00000_0000_00_010001100010", -- load, gr0, P1BOMB1ACTIVE
 464 => b"00011_0000_01_000000000000", -- sub, gr0
 465 => b"00000_0000_00_000000000001", -- 1
 466 => b"00111_0000_01_000000000000", -- bne
 467 => b"00000_0000_00_000111011101", -- P1BOMB2
 468 => b"00000_0000_00_010001100001", -- load, gr0, P1BOMB1TIME
 469 => b"00011_0000_01_000000000000", -- sub, gr0
 470 => b"00000_0000_00_000000000001", -- 1
 471 => b"00001_0000_10_010001100001", -- store, gr0, P1BOMB1TIME
 472 => b"00000_0000_01_000000000000", -- load, gr0
 473 => b"00000_0000_00_000000000000", -- 0
 474 => b"00011_0000_00_010001100001", -- sub, gr0, P1BOMB1TIME
 475 => b"00110_0000_01_000000000000", -- beq
 476 => b"00000_0000_00_001000100101", -- P1EXPLOSION1INIT
 477 => b"00000_0000_00_010001101000", -- load, gr0, P1BOMB2ACTIVE
 478 => b"00011_0000_01_000000000000", -- sub, gr0
 479 => b"00000_0000_00_000000000001", -- 1
 480 => b"00111_0000_01_000000000000", -- bne
 481 => b"00000_0000_00_000111101011", -- P1BOMB3
 482 => b"00000_0000_00_010001100111", -- load, gr0, P1BOMB2TIME
 483 => b"00011_0000_01_000000000000", -- sub, gr0
 484 => b"00000_0000_00_000000000001", -- 1
 485 => b"00001_0000_10_010001100111", -- store, gr0, P1BOMB2TIME
 486 => b"00000_0000_01_000000000000", -- load, gr0
 487 => b"00000_0000_00_000000000000", -- 0
 488 => b"00011_0000_00_010001100111", -- sub, gr0, P1BOMB2TIME
 489 => b"00110_0000_01_000000000000", -- beq
 490 => b"00000_0000_00_001000110111", -- P1EXPLOSION2INIT
 491 => b"00000_0000_00_010001101110", -- load, gr0, P1BOMB3ACTIVE
 492 => b"00011_0000_01_000000000000", -- sub, gr0
 493 => b"00000_0000_00_000000000001", -- 1
 494 => b"00111_0000_01_000000000000", -- bne
 495 => b"00000_0000_00_000111111001", -- P2BOMB1
 496 => b"00000_0000_00_010001101101", -- load, gr0, P1BOMB3TIME
 497 => b"00011_0000_01_000000000000", -- sub, gr0
 498 => b"00000_0000_00_000000000001", -- 1
 499 => b"00001_0000_10_010001101101", -- store, gr0, P1BOMB3TIME
 500 => b"00000_0000_01_000000000000", -- load, gr0
 501 => b"00000_0000_00_000000000000", -- 0
 502 => b"00011_0000_00_010001101101", -- sub, gr0, P1BOMB3TIME
 503 => b"00110_0000_01_000000000000", -- beq
 504 => b"00000_0000_00_001001001001", -- P1EXPLOSION3INIT
 505 => b"00000_0000_00_010001110100", -- load, gr0, P2BOMB1ACTIVE
 506 => b"00011_0000_01_000000000000", -- sub, gr0
 507 => b"00000_0000_00_000000000001", -- 1
 508 => b"00111_0000_01_000000000000", -- bne
 509 => b"00000_0000_00_001000000111", -- P2BOMB2
 510 => b"00000_0000_00_010001110011", -- load, gr0, P2BOMB1TIME
 511 => b"00011_0000_01_000000000000", -- sub, gr0
 512 => b"00000_0000_00_000000000001", -- 1
 513 => b"00001_0000_10_010001110011", -- store, gr0, P2BOMB1TIME
 514 => b"00000_0000_01_000000000000", -- load, gr0
 515 => b"00000_0000_00_000000000000", -- 0
 516 => b"00011_0000_00_010001110011", -- sub, gr0, P2BOMB1TIME
 517 => b"00110_0000_01_000000000000", -- beq
 518 => b"00000_0000_00_001001011011", -- P2EXPLOSION1INIT
 519 => b"00000_0000_00_010001111010", -- load, gr0, P2BOMB2ACTIVE
 520 => b"00011_0000_01_000000000000", -- sub, gr0
 521 => b"00000_0000_00_000000000001", -- 1
 522 => b"00111_0000_01_000000000000", -- bne
 523 => b"00000_0000_00_001000010101", -- P2BOMB3
 524 => b"00000_0000_00_010001111001", -- load, gr0, P2BOMB2TIME
 525 => b"00011_0000_01_000000000000", -- sub, gr0
 526 => b"00000_0000_00_000000000001", -- 1
 527 => b"00001_0000_10_010001111001", -- store, gr0, P2BOMB2TIME
 528 => b"00000_0000_01_000000000000", -- load, gr0
 529 => b"00000_0000_00_000000000000", -- 0
 530 => b"00011_0000_00_010001111001", -- sub, gr0, P2BOMB2TIME
 531 => b"00110_0000_01_000000000000", -- beq
 532 => b"00000_0000_00_001001101101", -- P2EXPLOSION2INIT
 533 => b"00000_0000_00_010010000000", -- load, gr0, P2BOMB3ACTIVE
 534 => b"00011_0000_01_000000000000", -- sub, gr0
 535 => b"00000_0000_00_000000000001", -- 1
 536 => b"00111_0000_01_000000000000", -- bne
 537 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 538 => b"00000_0000_00_010001111111", -- load, gr0, P2BOMB3TIME
 539 => b"00011_0000_01_000000000000", -- sub, gr0
 540 => b"00000_0000_00_000000000001", -- 1
 541 => b"00001_0000_10_010001111111", -- store, gr0, P2BOMB3TIME
 542 => b"00000_0000_01_000000000000", -- load, gr0
 543 => b"00000_0000_00_000000000000", -- 0
 544 => b"00011_0000_00_010001111111", -- sub, gr0, P2BOMB3TIME
 545 => b"00110_0000_01_000000000000", -- beq
 546 => b"00000_0000_00_001001111111", -- P2EXPLOSION3INIT
 547 => b"00100_0000_01_000000000000", -- jump
 548 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 549 => b"00000_0000_01_000000000000", -- load, gr0
 550 => b"00000_0000_00_000000000000", -- 0
 551 => b"00001_0000_10_010001100010", -- store, gr0, P1BOMB1ACTIVE
 552 => b"00000_0000_00_010001100000", -- load, gr0, P1BOMB1POS
 553 => b"00001_0000_10_010001100101", -- store, gr0, P1EXPLOSION1POS
 554 => b"00000_0000_01_000000000000", -- load, gr0
 555 => b"00000_0000_00_000000000001", -- 1
 556 => b"00001_0000_10_010001100100", -- store, gr0, P1EXPLOSION1ACTIVE
 557 => b"00000_0000_01_000000000000", -- load, gr0
 558 => b"00000_0000_00_000000000010", -- 2
 559 => b"00001_0000_10_010001100011", -- store, gr0, P1EXPLOSION1TIME
 560 => b"00000_0000_00_010010000100", -- load, gr0, P1BOMBCOUNT
 561 => b"00011_0000_01_000000000000", -- sub, gr0
 562 => b"00000_0000_00_000000000001", -- 1
 563 => b"00001_0000_10_010010000100", -- store, gr0, P1BOMBCOUNT
 564 => b"00000_0100_00_010001100000", -- load, gr4, P1BOMB1POS
 565 => b"00100_0000_01_000000000000", -- jump
 566 => b"00000_0000_00_001010010001", -- EXPLODE
 567 => b"00000_0000_01_000000000000", -- load, gr0
 568 => b"00000_0000_00_000000000000", -- 0
 569 => b"00001_0000_10_010001101000", -- store, gr0, P1BOMB2ACTIVE
 570 => b"00000_0000_00_010001100110", -- load, gr0, P1BOMB2POS
 571 => b"00001_0000_10_010001101011", -- store, gr0, P1EXPLOSION2POS
 572 => b"00000_0000_01_000000000000", -- load, gr0
 573 => b"00000_0000_00_000000000001", -- 1
 574 => b"00001_0000_10_010001101010", -- store, gr0, P1EXPLOSION2ACTIVE
 575 => b"00000_0000_01_000000000000", -- load, gr0
 576 => b"00000_0000_00_000000000010", -- 2
 577 => b"00001_0000_10_010001101001", -- store, gr0, P1EXPLOSION2TIME
 578 => b"00000_0000_00_010010000100", -- load, gr0, P1BOMBCOUNT
 579 => b"00011_0000_01_000000000000", -- sub, gr0
 580 => b"00000_0000_00_000000000001", -- 1
 581 => b"00001_0000_10_010010000100", -- store, gr0, P1BOMBCOUNT
 582 => b"00000_0100_00_010001100110", -- load, gr4, P1BOMB2POS
 583 => b"00100_0000_01_000000000000", -- jump
 584 => b"00000_0000_00_001010010001", -- EXPLODE
 585 => b"00000_0000_01_000000000000", -- load, gr0
 586 => b"00000_0000_00_000000000000", -- 0
 587 => b"00001_0000_10_010001101110", -- store, gr0, P1BOMB3ACTIVE
 588 => b"00000_0000_00_010001101100", -- load, gr0, P1BOMB3POS
 589 => b"00001_0000_10_010001110001", -- store, gr0, P1EXPLOSION3POS
 590 => b"00000_0000_01_000000000000", -- load, gr0
 591 => b"00000_0000_00_000000000001", -- 1
 592 => b"00001_0000_10_010001110000", -- store, gr0, P1EXPLOSION3ACTIVE
 593 => b"00000_0000_01_000000000000", -- load, gr0
 594 => b"00000_0000_00_000000000010", -- 2
 595 => b"00001_0000_10_010001101111", -- store, gr0, P1EXPLOSION3TIME
 596 => b"00000_0000_00_010010000100", -- load, gr0, P1BOMBCOUNT
 597 => b"00011_0000_01_000000000000", -- sub, gr0
 598 => b"00000_0000_00_000000000001", -- 1
 599 => b"00001_0000_10_010010000100", -- store, gr0, P1BOMBCOUNT
 600 => b"00000_0100_00_010001101100", -- load, gr4, P1BOMB3POS
 601 => b"00100_0000_01_000000000000", -- jump
 602 => b"00000_0000_00_001010010001", -- EXPLODE
 603 => b"00000_0000_01_000000000000", -- load, gr0
 604 => b"00000_0000_00_000000000000", -- 0
 605 => b"00001_0000_10_010001110100", -- store, gr0, P2BOMB1ACTIVE
 606 => b"00000_0000_00_010001110010", -- load, gr0, P2BOMB1POS
 607 => b"00001_0000_10_010001110111", -- store, gr0, P2EXPLOSION1POS
 608 => b"00000_0000_01_000000000000", -- load, gr0
 609 => b"00000_0000_00_000000000001", -- 1
 610 => b"00001_0000_10_010001110110", -- store, gr0, P2EXPLOSION1ACTIVE
 611 => b"00000_0000_01_000000000000", -- load, gr0
 612 => b"00000_0000_00_000000000010", -- 2
 613 => b"00001_0000_10_010001110101", -- store, gr0, P2EXPLOSION1TIME
 614 => b"00000_0000_00_010010000101", -- load, gr0, P2BOMBCOUNT
 615 => b"00011_0000_01_000000000000", -- sub, gr0
 616 => b"00000_0000_00_000000000001", -- 1
 617 => b"00001_0000_10_010010000101", -- store, gr0, P2BOMBCOUNT
 618 => b"00000_0100_00_010001110010", -- load, gr4, P2BOMB1POS
 619 => b"00100_0000_01_000000000000", -- jump
 620 => b"00000_0000_00_001010010001", -- EXPLODE
 621 => b"00000_0000_01_000000000000", -- load, gr0
 622 => b"00000_0000_00_000000000000", -- 0
 623 => b"00001_0000_10_010001111010", -- store, gr0, P2BOMB2ACTIVE
 624 => b"00000_0000_00_010001111000", -- load, gr0, P2BOMB2POS
 625 => b"00001_0000_10_010001111101", -- store, gr0, P2EXPLOSION2POS
 626 => b"00000_0000_01_000000000000", -- load, gr0
 627 => b"00000_0000_00_000000000001", -- 1
 628 => b"00001_0000_10_010001111100", -- store, gr0, P2EXPLOSION2ACTIVE
 629 => b"00000_0000_01_000000000000", -- load, gr0
 630 => b"00000_0000_00_000000000010", -- 2
 631 => b"00001_0000_10_010001111011", -- store, gr0, P2EXPLOSION2TIME
 632 => b"00000_0000_00_010010000101", -- load, gr0, P2BOMBCOUNT
 633 => b"00011_0000_01_000000000000", -- sub, gr0
 634 => b"00000_0000_00_000000000001", -- 1
 635 => b"00001_0000_10_010010000101", -- store, gr0, P2BOMBCOUNT
 636 => b"00000_0100_00_010001111000", -- load, gr4, P2BOMB2POS
 637 => b"00100_0000_01_000000000000", -- jump
 638 => b"00000_0000_00_001010010001", -- EXPLODE
 639 => b"00000_0000_01_000000000000", -- load, gr0
 640 => b"00000_0000_00_000000000000", -- 0
 641 => b"00001_0000_10_010010000000", -- store, gr0, P2BOMB3ACTIVE
 642 => b"00000_0000_00_010001111110", -- load, gr0, P2BOMB3POS
 643 => b"00001_0000_10_010010000011", -- store, gr0, P2EXPLOSION3POS
 644 => b"00000_0000_01_000000000000", -- load, gr0
 645 => b"00000_0000_00_000000000001", -- 1
 646 => b"00001_0000_10_010010000010", -- store, gr0, P2EXPLOSION3ACTIVE
 647 => b"00000_0000_01_000000000000", -- load, gr0
 648 => b"00000_0000_00_000000000010", -- 2
 649 => b"00001_0000_10_010010000001", -- store, gr0, P2EXPLOSION3TIME
 650 => b"00000_0000_00_010010000101", -- load, gr0, P2BOMBCOUNT
 651 => b"00011_0000_01_000000000000", -- sub, gr0
 652 => b"00000_0000_00_000000000001", -- 1
 653 => b"00001_0000_10_010010000101", -- store, gr0, P2BOMBCOUNT
 654 => b"00000_0100_00_010001111110", -- load, gr4, P2BOMB3POS
 655 => b"00100_0000_01_000000000000", -- jump
 656 => b"00000_0000_00_001010010001", -- EXPLODE
 657 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 658 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 659 => b"00000_0011_00_010010010001", -- load, gr3, EXPLOSION
 660 => b"10000_0010_00_000000000000", -- tpoint, gr2
 661 => b"01110_0011_00_000000000000", -- twrite, gr3
 662 => b"00010_0010_01_000000000000", -- add, gr2
 663 => b"00000_0000_00_000000000001", -- 1
 664 => b"10000_0010_00_000000000000", -- tpoint, gr2
 665 => b"01111_0000_00_000000000000", -- tread, gr0
 666 => b"00001_0000_10_010010001011", -- store, gr0, MOVE
 667 => b"00000_0111_00_010010001011", -- load, gr7, MOVE
 668 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 669 => b"00110_0000_01_000000000000", -- beq
 670 => b"00000_0000_00_001010101011", -- EXPLODELEFT
 671 => b"01110_0011_00_000000000000", -- twrite, gr3
 672 => b"00011_0111_00_010010010000", -- sub, gr7, BREAKABLE
 673 => b"00110_0000_01_000000000000", -- beq
 674 => b"00000_0000_00_001010101011", -- EXPLODELEFT
 675 => b"00010_0010_01_000000000000", -- add, gr2
 676 => b"00000_0000_00_000000000001", -- 1
 677 => b"10000_0010_00_000000000000", -- tpoint, gr2
 678 => b"01111_0000_00_000000000000", -- tread, gr0
 679 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 680 => b"00110_0000_01_000000000000", -- beq
 681 => b"00000_0000_00_001010101011", -- EXPLODELEFT
 682 => b"01110_0011_00_000000000000", -- twrite, gr3
 683 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 684 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 685 => b"00011_0010_01_000000000000", -- sub, gr2
 686 => b"00000_0000_00_000000000001", -- 1
 687 => b"10000_0010_00_000000000000", -- tpoint, gr2
 688 => b"01111_0000_00_000000000000", -- tread, gr0
 689 => b"00001_0000_10_010010001011", -- store, gr0, MOVE
 690 => b"00000_0111_00_010010001011", -- load, gr7, MOVE
 691 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 692 => b"00110_0000_01_000000000000", -- beq
 693 => b"00000_0000_00_001011000010", -- EXPLODEDOWN
 694 => b"01110_0011_00_000000000000", -- twrite, gr3
 695 => b"00011_0111_00_010010010000", -- sub, gr7, BREAKABLE
 696 => b"00110_0000_01_000000000000", -- beq
 697 => b"00000_0000_00_001011000010", -- EXPLODEDOWN
 698 => b"00011_0010_01_000000000000", -- sub, gr2
 699 => b"00000_0000_00_000000000001", -- 1
 700 => b"10000_0010_00_000000000000", -- tpoint, gr2
 701 => b"01111_0000_00_000000000000", -- tread, gr0
 702 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 703 => b"00110_0000_01_000000000000", -- beq
 704 => b"00000_0000_00_001011000010", -- EXPLODEDOWN
 705 => b"01110_0011_00_000000000000", -- twrite, gr3
 706 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 707 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 708 => b"00010_0010_01_000000000000", -- add, gr2
 709 => b"00000_0000_00_000000001111", -- 15
 710 => b"10000_0010_00_000000000000", -- tpoint, gr2
 711 => b"01111_0000_00_000000000000", -- tread, gr0
 712 => b"00001_0000_10_010010001011", -- store, gr0, MOVE
 713 => b"00000_0111_00_010010001011", -- load, gr7, MOVE
 714 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 715 => b"00110_0000_01_000000000000", -- beq
 716 => b"00000_0000_00_001011011001", -- EXPLODEUP
 717 => b"01110_0011_00_000000000000", -- twrite, gr3
 718 => b"00011_0111_00_010010010000", -- sub, gr7, BREAKABLE
 719 => b"00110_0000_01_000000000000", -- beq
 720 => b"00000_0000_00_001011011001", -- EXPLODEUP
 721 => b"00010_0010_01_000000000000", -- add, gr2
 722 => b"00000_0000_00_000000001111", -- 15
 723 => b"10000_0010_00_000000000000", -- tpoint, gr2
 724 => b"01111_0000_00_000000000000", -- tread, gr0
 725 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 726 => b"00110_0000_01_000000000000", -- beq
 727 => b"00000_0000_00_001011011001", -- EXPLODEUP
 728 => b"01110_0011_00_000000000000", -- twrite, gr3
 729 => b"00001_0100_10_010010001011", -- store, gr4, MOVE
 730 => b"00000_0010_00_010010001011", -- load, gr2, MOVE
 731 => b"00011_0010_01_000000000000", -- sub, gr2
 732 => b"00000_0000_00_000000001111", -- 15
 733 => b"10000_0010_00_000000000000", -- tpoint, gr2
 734 => b"01111_0000_00_000000000000", -- tread, gr0
 735 => b"00001_0000_10_010010001011", -- store, gr0, MOVE
 736 => b"00000_0111_00_010010001011", -- load, gr7, MOVE
 737 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 738 => b"00110_0000_01_000000000000", -- beq
 739 => b"00000_0000_00_000111001111", -- TICKBOMBS
 740 => b"01110_0011_00_000000000000", -- twrite, gr3
 741 => b"00011_0111_00_010010010000", -- sub, gr7, BREAKABLE
 742 => b"00110_0000_01_000000000000", -- beq
 743 => b"00000_0000_00_000111001111", -- TICKBOMBS
 744 => b"00011_0010_01_000000000000", -- sub, gr2
 745 => b"00000_0000_00_000000001111", -- 15
 746 => b"10000_0010_00_000000000000", -- tpoint, gr2
 747 => b"01111_0000_00_000000000000", -- tread, gr0
 748 => b"00011_0000_00_010010001111", -- sub, gr0, WALL
 749 => b"00110_0000_01_000000000000", -- beq
 750 => b"00000_0000_00_000111001111", -- TICKBOMBS
 751 => b"01110_0011_00_000000000000", -- twrite, gr3
 752 => b"00100_0000_01_000000000000", -- jump
 753 => b"00000_0000_00_000111001111", -- TICKBOMBS
 754 => b"10101_0000_01_000000000000", -- btn1
 755 => b"00000_0000_00_001011111000", -- BTN1
 756 => b"11010_0000_01_000000000000", -- btn2
 757 => b"00000_0000_00_001101011001", -- BTN2
 758 => b"00100_0000_01_000000000000", -- jump
 759 => b"00000_0000_00_000001101000", -- BUTTON_R
 760 => b"00000_0000_00_010001011100", -- load, gr0, P1DEAD
 761 => b"00011_0000_01_000000000000", -- sub, gr0
 762 => b"00000_0000_00_000000000001", -- 1
 763 => b"00110_0000_01_000000000000", -- beq
 764 => b"00000_0000_00_000000000000", -- INIT
 765 => b"00000_0000_00_010010000100", -- load, gr0, P1BOMBCOUNT
 766 => b"00011_0000_00_010010000110", -- sub, gr0, MAXBOMBS
 767 => b"00110_0000_01_000000000000", -- beq
 768 => b"00000_0000_00_001011110100", -- BTN1_R
 769 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 770 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 771 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
 772 => b"01000_0000_01_000000000000", -- mul, gr0
 773 => b"00000_0000_00_000000001111", -- 15
 774 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
 775 => b"10000_0000_00_000000000000", -- tpoint, gr0
 776 => b"01111_0001_00_000000000000", -- tread, gr1
 777 => b"00011_0001_00_010010010010", -- sub, gr1, EGG
 778 => b"00110_0000_01_000000000000", -- beq
 779 => b"00000_0000_00_001011110100", -- BTN1_R
 780 => b"00000_0000_00_010001100010", -- load, gr0, P1BOMB1ACTIVE
 781 => b"00011_0000_01_000000000000", -- sub, gr0
 782 => b"00000_0000_00_000000000000", -- 0
 783 => b"00110_0000_01_000000000000", -- beq
 784 => b"00000_0000_00_001100100011", -- P1PLACEBOMB1
 785 => b"00000_0000_00_010001101000", -- load, gr0, P1BOMB2ACTIVE
 786 => b"00011_0000_01_000000000000", -- sub, gr0
 787 => b"00000_0000_00_000000000000", -- 0
 788 => b"00110_0000_01_000000000000", -- beq
 789 => b"00000_0000_00_001100110101", -- P1PLACEBOMB2
 790 => b"00000_0000_00_010001101110", -- load, gr0, P1BOMB3ACTIVE
 791 => b"00011_0000_01_000000000000", -- sub, gr0
 792 => b"00000_0000_00_000000000000", -- 0
 793 => b"00110_0000_01_000000000000", -- beq
 794 => b"00000_0000_00_001101000111", -- P1PLACEBOMB3
 795 => b"00100_0000_01_000000000000", -- jump
 796 => b"00000_0000_00_001011110100", -- BTN1_R
 797 => b"00000_0000_00_010010000100", -- load, gr0, P1BOMBCOUNT
 798 => b"00010_0000_01_000000000000", -- add, gr0
 799 => b"00000_0000_00_000000000001", -- 1
 800 => b"00001_0000_10_010010000100", -- store, gr0, P1BOMBCOUNT
 801 => b"00100_0000_01_000000000000", -- jump
 802 => b"00000_0000_00_001011110100", -- BTN1_R
 803 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 804 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 805 => b"00000_0011_00_010010001000", -- load, gr3, YPOS1
 806 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 807 => b"01000_0011_01_000000000000", -- mul, gr3
 808 => b"00000_0000_00_000000001111", -- 15
 809 => b"00010_0011_00_010010000111", -- add, gr3, XPOS1
 810 => b"10000_0011_00_000000000000", -- tpoint, gr3
 811 => b"01110_0010_00_000000000000", -- twrite, gr2
 812 => b"00000_0000_01_000000000000", -- load, gr0
 813 => b"00000_0000_00_000000000001", -- 1
 814 => b"00001_0000_10_010001100010", -- store, gr0, P1BOMB1ACTIVE
 815 => b"00001_0011_10_010001100000", -- store, gr3, P1BOMB1POS
 816 => b"00000_0000_01_000000000000", -- load, gr0
 817 => b"00000_0000_00_000000010000", -- 16
 818 => b"00001_0000_10_010001100001", -- store, gr0, P1BOMB1TIME
 819 => b"00100_0000_01_000000000000", -- jump
 820 => b"00000_0000_00_001100011101", -- P1INCREASEBOMBCOUNTER
 821 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 822 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 823 => b"00000_0011_00_010010001000", -- load, gr3, YPOS1
 824 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 825 => b"01000_0011_01_000000000000", -- mul, gr3
 826 => b"00000_0000_00_000000001111", -- 15
 827 => b"00010_0011_00_010010000111", -- add, gr3, XPOS1
 828 => b"10000_0011_00_000000000000", -- tpoint, gr3
 829 => b"01110_0010_00_000000000000", -- twrite, gr2
 830 => b"00000_0000_01_000000000000", -- load, gr0
 831 => b"00000_0000_00_000000000001", -- 1
 832 => b"00001_0000_10_010001101000", -- store, gr0, P1BOMB2ACTIVE
 833 => b"00001_0011_10_010001100110", -- store, gr3, P1BOMB2POS
 834 => b"00000_0000_01_000000000000", -- load, gr0
 835 => b"00000_0000_00_000000010000", -- 16
 836 => b"00001_0000_10_010001100111", -- store, gr0, P1BOMB2TIME
 837 => b"00100_0000_01_000000000000", -- jump
 838 => b"00000_0000_00_001100011101", -- P1INCREASEBOMBCOUNTER
 839 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 840 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 841 => b"00000_0011_00_010010001000", -- load, gr3, YPOS1
 842 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 843 => b"01000_0011_01_000000000000", -- mul, gr3
 844 => b"00000_0000_00_000000001111", -- 15
 845 => b"00010_0011_00_010010000111", -- add, gr3, XPOS1
 846 => b"10000_0011_00_000000000000", -- tpoint, gr3
 847 => b"01110_0010_00_000000000000", -- twrite, gr2
 848 => b"00000_0000_01_000000000000", -- load, gr0
 849 => b"00000_0000_00_000000000001", -- 1
 850 => b"00001_0000_10_010001101110", -- store, gr0, P1BOMB3ACTIVE
 851 => b"00001_0011_10_010001101100", -- store, gr3, P1BOMB3POS
 852 => b"00000_0000_01_000000000000", -- load, gr0
 853 => b"00000_0000_00_000000010000", -- 16
 854 => b"00001_0000_10_010001101101", -- store, gr0, P1BOMB3TIME
 855 => b"00100_0000_01_000000000000", -- jump
 856 => b"00000_0000_00_001100011101", -- P1INCREASEBOMBCOUNTER
 857 => b"00000_0000_00_010001011101", -- load, gr0, P2DEAD
 858 => b"00011_0000_01_000000000000", -- sub, gr0
 859 => b"00000_0000_00_000000000001", -- 1
 860 => b"00110_0000_01_000000000000", -- beq
 861 => b"00000_0000_00_000000000000", -- INIT
 862 => b"00000_0000_00_010010000101", -- load, gr0, P2BOMBCOUNT
 863 => b"00011_0000_00_010010000110", -- sub, gr0, MAXBOMBS
 864 => b"00110_0000_01_000000000000", -- beq
 865 => b"00000_0000_00_001011110110", -- BTN2_R
 866 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 867 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 868 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
 869 => b"01000_0000_01_000000000000", -- mul, gr0
 870 => b"00000_0000_00_000000001111", -- 15
 871 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
 872 => b"10000_0000_00_000000000000", -- tpoint, gr0
 873 => b"01111_0001_00_000000000000", -- tread, gr1
 874 => b"00011_0001_00_010010010010", -- sub, gr1, EGG
 875 => b"00110_0000_01_000000000000", -- beq
 876 => b"00000_0000_00_001011110110", -- BTN2_R
 877 => b"00000_0000_00_010001110100", -- load, gr0, P2BOMB1ACTIVE
 878 => b"00011_0000_01_000000000000", -- sub, gr0
 879 => b"00000_0000_00_000000000000", -- 0
 880 => b"00110_0000_01_000000000000", -- beq
 881 => b"00000_0000_00_001110000010", -- P2PLACEBOMB1
 882 => b"00000_0000_00_010001111010", -- load, gr0, P2BOMB2ACTIVE
 883 => b"00011_0000_01_000000000000", -- sub, gr0
 884 => b"00000_0000_00_000000000000", -- 0
 885 => b"00110_0000_01_000000000000", -- beq
 886 => b"00000_0000_00_001110010100", -- P2PLACEBOMB2
 887 => b"00000_0000_00_010010000000", -- load, gr0, P2BOMB3ACTIVE
 888 => b"00011_0000_01_000000000000", -- sub, gr0
 889 => b"00000_0000_00_000000000000", -- 0
 890 => b"00110_0000_01_000000000000", -- beq
 891 => b"00000_0000_00_001110100110", -- P2PLACEBOMB3
 892 => b"00000_0000_00_010010000101", -- load, gr0, P2BOMBCOUNT
 893 => b"00010_0000_01_000000000000", -- add, gr0
 894 => b"00000_0000_00_000000000001", -- 1
 895 => b"00001_0000_10_010010000101", -- store, gr0, P2BOMBCOUNT
 896 => b"00100_0000_01_000000000000", -- jump
 897 => b"00000_0000_00_001011110110", -- BTN2_R
 898 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 899 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 900 => b"00000_0011_00_010010001010", -- load, gr3, YPOS2
 901 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 902 => b"01000_0011_01_000000000000", -- mul, gr3
 903 => b"00000_0000_00_000000001111", -- 15
 904 => b"00010_0011_00_010010001001", -- add, gr3, XPOS2
 905 => b"10000_0011_00_000000000000", -- tpoint, gr3
 906 => b"01110_0010_00_000000000000", -- twrite, gr2
 907 => b"00000_0000_01_000000000000", -- load, gr0
 908 => b"00000_0000_00_000000000001", -- 1
 909 => b"00001_0000_10_010001110100", -- store, gr0, P2BOMB1ACTIVE
 910 => b"00001_0011_10_010001110010", -- store, gr3, P2BOMB1POS
 911 => b"00000_0000_01_000000000000", -- load, gr0
 912 => b"00000_0000_00_000000010000", -- 16
 913 => b"00001_0000_10_010001110011", -- store, gr0, P2BOMB1TIME
 914 => b"00100_0000_01_000000000000", -- jump
 915 => b"00000_0000_00_001101111100", -- P2INCREASEBOMBCOUNTER
 916 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 917 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 918 => b"00000_0011_00_010010001010", -- load, gr3, YPOS2
 919 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 920 => b"01000_0011_01_000000000000", -- mul, gr3
 921 => b"00000_0000_00_000000001111", -- 15
 922 => b"00010_0011_00_010010001001", -- add, gr3, XPOS2
 923 => b"10000_0011_00_000000000000", -- tpoint, gr3
 924 => b"01110_0010_00_000000000000", -- twrite, gr2
 925 => b"00000_0000_01_000000000000", -- load, gr0
 926 => b"00000_0000_00_000000000001", -- 1
 927 => b"00001_0000_10_010001111010", -- store, gr0, P2BOMB2ACTIVE
 928 => b"00001_0011_10_010001111000", -- store, gr3, P2BOMB2POS
 929 => b"00000_0000_01_000000000000", -- load, gr0
 930 => b"00000_0000_00_000000010000", -- 16
 931 => b"00001_0000_10_010001111001", -- store, gr0, P2BOMB2TIME
 932 => b"00100_0000_01_000000000000", -- jump
 933 => b"00000_0000_00_001101111100", -- P2INCREASEBOMBCOUNTER
 934 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
 935 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
 936 => b"00000_0011_00_010010001010", -- load, gr3, YPOS2
 937 => b"00000_0010_00_010010010010", -- load, gr2, EGG
 938 => b"01000_0011_01_000000000000", -- mul, gr3
 939 => b"00000_0000_00_000000001111", -- 15
 940 => b"00010_0011_00_010010001001", -- add, gr3, XPOS2
 941 => b"10000_0011_00_000000000000", -- tpoint, gr3
 942 => b"01110_0010_00_000000000000", -- twrite, gr2
 943 => b"00000_0000_01_000000000000", -- load, gr0
 944 => b"00000_0000_00_000000000001", -- 1
 945 => b"00001_0000_10_010010000000", -- store, gr0, P2BOMB3ACTIVE
 946 => b"00001_0011_10_010001111110", -- store, gr3, P2BOMB3POS
 947 => b"00000_0000_01_000000000000", -- load, gr0
 948 => b"00000_0000_00_000000010000", -- 16
 949 => b"00001_0000_10_010001111111", -- store, gr0, P2BOMB3TIME
 950 => b"00100_0000_01_000000000000", -- jump
 951 => b"00000_0000_00_001101111100", -- P2INCREASEBOMBCOUNTER
 952 => b"00000_0000_00_010001011100", -- load, gr0, P1DEAD
 953 => b"00011_0000_01_000000000000", -- sub, gr0
 954 => b"00000_0000_00_000000000001", -- 1
 955 => b"00110_0000_01_000000000000", -- beq
 956 => b"00000_0000_00_001111000101", -- J2
 957 => b"10001_0000_01_000000000000", -- joy1r
 958 => b"00000_0000_00_001111010100", -- P1R
 959 => b"10011_0000_01_000000000000", -- joy1l
 960 => b"00000_0000_00_001111110110", -- P1L
 961 => b"10010_0000_01_000000000000", -- joy1u
 962 => b"00000_0000_00_001111100101", -- P1U
 963 => b"10100_0000_01_000000000000", -- joy1d
 964 => b"00000_0000_00_010000000111", -- P1D
 965 => b"00000_0000_00_010001011101", -- load, gr0, P2DEAD
 966 => b"00011_0000_01_000000000000", -- sub, gr0
 967 => b"00000_0000_00_000000000001", -- 1
 968 => b"00110_0000_01_000000000000", -- beq
 969 => b"00000_0000_00_000001100110", -- CONTROL_R
 970 => b"10110_0000_01_000000000000", -- joy2r
 971 => b"00000_0000_00_010000011000", -- P2R
 972 => b"11000_0000_01_000000000000", -- joy2l
 973 => b"00000_0000_00_010000111010", -- P2L
 974 => b"10111_0000_01_000000000000", -- joy2u
 975 => b"00000_0000_00_010000101001", -- P2U
 976 => b"11001_0000_01_000000000000", -- joy2d
 977 => b"00000_0000_00_010001001011", -- P2D
 978 => b"00100_0000_01_000000000000", -- jump
 979 => b"00000_0000_00_000001100110", -- CONTROL_R
 980 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 981 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 982 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
 983 => b"01000_0000_01_000000000000", -- mul, gr0
 984 => b"00000_0000_00_000000001111", -- 15
 985 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
 986 => b"00010_0000_01_000000000000", -- add, gr0
 987 => b"00000_0000_00_000000000001", -- 1
 988 => b"10000_0000_00_000000000000", -- tpoint, gr0
 989 => b"01111_0001_00_000000000000", -- tread, gr1
 990 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
 991 => b"00111_0000_01_000000000000", -- bne
 992 => b"00000_0000_00_001111000001", -- J1
 993 => b"00010_1100_01_000000000000", -- add, gr12
 994 => b"00000_0000_00_000000000001", -- 1
 995 => b"00100_0000_01_000000000000", -- jump
 996 => b"00000_0000_00_001111000001", -- J1
 997 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
 998 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
 999 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
1000 => b"00011_0000_01_000000000000", -- sub, gr0
1001 => b"00000_0000_00_000000000001", -- 1
1002 => b"01000_0000_01_000000000000", -- mul, gr0
1003 => b"00000_0000_00_000000001111", -- 15
1004 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
1005 => b"10000_0000_00_000000000000", -- tpoint, gr0
1006 => b"01111_0001_00_000000000000", -- tread, gr1
1007 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1008 => b"00111_0000_01_000000000000", -- bne
1009 => b"00000_0000_00_001111000101", -- J2
1010 => b"00011_1101_01_000000000000", -- sub, gr13
1011 => b"00000_0000_00_000000000001", -- 1
1012 => b"00100_0000_01_000000000000", -- jump
1013 => b"00000_0000_00_001111000101", -- J2
1014 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
1015 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
1016 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
1017 => b"01000_0000_01_000000000000", -- mul, gr0
1018 => b"00000_0000_00_000000001111", -- 15
1019 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
1020 => b"00011_0000_01_000000000000", -- sub, gr0
1021 => b"00000_0000_00_000000000001", -- 1
1022 => b"10000_0000_00_000000000000", -- tpoint, gr0
1023 => b"01111_0001_00_000000000000", -- tread, gr1
1024 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1025 => b"00111_0000_01_000000000000", -- bne
1026 => b"00000_0000_00_001111000001", -- J1
1027 => b"00011_1100_01_000000000000", -- sub, gr12
1028 => b"00000_0000_00_000000000001", -- 1
1029 => b"00100_0000_01_000000000000", -- jump
1030 => b"00000_0000_00_001111000001", -- J1
1031 => b"00001_1100_10_010010000111", -- store, gr12, XPOS1
1032 => b"00001_1101_10_010010001000", -- store, gr13, YPOS1
1033 => b"00000_0000_00_010010001000", -- load, gr0, YPOS1
1034 => b"00010_0000_01_000000000000", -- add, gr0
1035 => b"00000_0000_00_000000000001", -- 1
1036 => b"01000_0000_01_000000000000", -- mul, gr0
1037 => b"00000_0000_00_000000001111", -- 15
1038 => b"00010_0000_00_010010000111", -- add, gr0, XPOS1
1039 => b"10000_0000_00_000000000000", -- tpoint, gr0
1040 => b"01111_0001_00_000000000000", -- tread, gr1
1041 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1042 => b"00111_0000_01_000000000000", -- bne
1043 => b"00000_0000_00_001111000101", -- J2
1044 => b"00010_1101_01_000000000000", -- add, gr13
1045 => b"00000_0000_00_000000000001", -- 1
1046 => b"00100_0000_01_000000000000", -- jump
1047 => b"00000_0000_00_001111000101", -- J2
1048 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
1049 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
1050 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
1051 => b"01000_0000_01_000000000000", -- mul, gr0
1052 => b"00000_0000_00_000000001111", -- 15
1053 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
1054 => b"00010_0000_01_000000000000", -- add, gr0
1055 => b"00000_0000_00_000000000001", -- 1
1056 => b"10000_0000_00_000000000000", -- tpoint, gr0
1057 => b"01111_0001_00_000000000000", -- tread, gr1
1058 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1059 => b"00111_0000_01_000000000000", -- bne
1060 => b"00000_0000_00_001111001110", -- J3
1061 => b"00010_1110_01_000000000000", -- add, gr14
1062 => b"00000_0000_00_000000000001", -- 1
1063 => b"00100_0000_01_000000000000", -- jump
1064 => b"00000_0000_00_001111001110", -- J3
1065 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
1066 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
1067 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
1068 => b"00011_0000_01_000000000000", -- sub, gr0
1069 => b"00000_0000_00_000000000001", -- 1
1070 => b"01000_0000_01_000000000000", -- mul, gr0
1071 => b"00000_0000_00_000000001111", -- 15
1072 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
1073 => b"10000_0000_00_000000000000", -- tpoint, gr0
1074 => b"01111_0001_00_000000000000", -- tread, gr1
1075 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1076 => b"00111_0000_01_000000000000", -- bne
1077 => b"00000_0000_00_000001100110", -- CONTROL_R
1078 => b"00011_1111_01_000000000000", -- sub, gr15
1079 => b"00000_0000_00_000000000001", -- 1
1080 => b"00100_0000_01_000000000000", -- jump
1081 => b"00000_0000_00_000001100110", -- CONTROL_R
1082 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
1083 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
1084 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
1085 => b"01000_0000_01_000000000000", -- mul, gr0
1086 => b"00000_0000_00_000000001111", -- 15
1087 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
1088 => b"00011_0000_01_000000000000", -- sub, gr0
1089 => b"00000_0000_00_000000000001", -- 1
1090 => b"10000_0000_00_000000000000", -- tpoint, gr0
1091 => b"01111_0001_00_000000000000", -- tread, gr1
1092 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1093 => b"00111_0000_01_000000000000", -- bne
1094 => b"00000_0000_00_001111001110", -- J3
1095 => b"00011_1110_01_000000000000", -- sub, gr14
1096 => b"00000_0000_00_000000000001", -- 1
1097 => b"00100_0000_01_000000000000", -- jump
1098 => b"00000_0000_00_001111001110", -- J3
1099 => b"00001_1110_10_010010001001", -- store, gr14, XPOS2
1100 => b"00001_1111_10_010010001010", -- store, gr15, YPOS2
1101 => b"00000_0000_00_010010001010", -- load, gr0, YPOS2
1102 => b"00010_0000_01_000000000000", -- add, gr0
1103 => b"00000_0000_00_000000000001", -- 1
1104 => b"01000_0000_01_000000000000", -- mul, gr0
1105 => b"00000_0000_00_000000001111", -- 15
1106 => b"00010_0000_00_010010001001", -- add, gr0, XPOS2
1107 => b"10000_0000_00_000000000000", -- tpoint, gr0
1108 => b"01111_0001_00_000000000000", -- tread, gr1
1109 => b"00011_0001_00_010010001110", -- sub, gr1, GRASS
1110 => b"00111_0000_01_000000000000", -- bne
1111 => b"00000_0000_00_000001100110", -- CONTROL_R
1112 => b"00010_1111_01_000000000000", -- add, gr15
1113 => b"00000_0000_00_000000000001", -- 1
1114 => b"00100_0000_01_000000000000", -- jump
1115 => b"00000_0000_00_000001100110", -- CONTROL_R
1116 => b"00000_0000_00_000000000000", -- 0
1117 => b"00000_0000_00_000000000000", -- 0
1118 => b"00000_0000_00_000000000000", -- 0
1119 => b"00000_0000_00_000000000000", -- 0
1120 => b"00000_0000_00_000000000000", -- 0
1121 => b"00000_0000_00_000000000000", -- 0
1122 => b"00000_0000_00_000000000000", -- 0
1123 => b"00000_0000_00_000000000000", -- 0
1124 => b"00000_0000_00_000000000000", -- 0
1125 => b"00000_0000_00_000000000000", -- 0
1126 => b"00000_0000_00_000000000000", -- 0
1127 => b"00000_0000_00_000000000000", -- 0
1128 => b"00000_0000_00_000000000000", -- 0
1129 => b"00000_0000_00_000000000000", -- 0
1130 => b"00000_0000_00_000000000000", -- 0
1131 => b"00000_0000_00_000000000000", -- 0
1132 => b"00000_0000_00_000000000000", -- 0
1133 => b"00000_0000_00_000000000000", -- 0
1134 => b"00000_0000_00_000000000000", -- 0
1135 => b"00000_0000_00_000000000000", -- 0
1136 => b"00000_0000_00_000000000000", -- 0
1137 => b"00000_0000_00_000000000000", -- 0
1138 => b"00000_0000_00_000000000000", -- 0
1139 => b"00000_0000_00_000000000000", -- 0
1140 => b"00000_0000_00_000000000000", -- 0
1141 => b"00000_0000_00_000000000000", -- 0
1142 => b"00000_0000_00_000000000000", -- 0
1143 => b"00000_0000_00_000000000000", -- 0
1144 => b"00000_0000_00_000000000000", -- 0
1145 => b"00000_0000_00_000000000000", -- 0
1146 => b"00000_0000_00_000000000000", -- 0
1147 => b"00000_0000_00_000000000000", -- 0
1148 => b"00000_0000_00_000000000000", -- 0
1149 => b"00000_0000_00_000000000000", -- 0
1150 => b"00000_0000_00_000000000000", -- 0
1151 => b"00000_0000_00_000000000000", -- 0
1152 => b"00000_0000_00_000000000000", -- 0
1153 => b"00000_0000_00_000000000000", -- 0
1154 => b"00000_0000_00_000000000000", -- 0
1155 => b"00000_0000_00_000000000000", -- 0
1156 => b"00000_0000_00_000000000000", -- 0
1157 => b"00000_0000_00_000000000000", -- 0
1158 => b"00000_0000_00_000000000011", -- 3
1159 => b"00000_0000_00_000000000000", -- 0
1160 => b"00000_0000_00_000000000000", -- 0
1161 => b"00000_0000_00_000000000000", -- 0
1162 => b"00000_0000_00_000000000000", -- 0
1163 => b"00000_0000_00_000000000000", -- 0
1164 => b"00000_0000_00_000000000000", -- 0
1165 => b"00000_0000_00_000000000000", -- 0
1166 => b"00000_0000_00_000000000000", -- 0
1167 => b"00000_0000_00_000000000001", -- 1
1168 => b"00000_0000_00_000000000010", -- 2
1169 => b"00000_0000_00_000000000011", -- 3
1170 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
