library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_001000000111", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000101001101", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011000100", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000010000", -- BOOM1
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000001101010", -- BOOM2
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  16 => b"00000_0000_00_001010101001", -- load, gr0, P1EXPLOSION1ACTIVE
  17 => b"00011_0000_01_000000000000", -- sub, gr0
  18 => b"00000_0000_00_000000000001", -- 1
  19 => b"00111_0000_01_000000000000", -- bne
  20 => b"00000_0000_00_000000001100", -- BOOM1_R
  21 => b"00000_0000_00_001010101000", -- load, gr0, P1EXPLOSION1TIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000001", -- 1
  24 => b"00001_0000_10_001010101000", -- store, gr0, P1EXPLOSION1TIME
  25 => b"00000_0000_00_001010101000", -- load, gr0, P1EXPLOSION1TIME
  26 => b"00011_0000_01_000000000000", -- sub, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00111_0000_01_000000000000", -- bne
  29 => b"00000_0000_00_000000001100", -- BOOM1_R
  30 => b"00000_0000_01_000000000000", -- load, gr0
  31 => b"00000_0000_00_000000000000", -- 0
  32 => b"00001_0000_10_001010101001", -- store, gr0, P1EXPLOSION1ACTIVE
  33 => b"00000_0010_00_001010101010", -- load, gr2, P1EXPLOSION1POS
  34 => b"00000_0011_00_001011010011", -- load, gr3, GRASS
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01110_0011_00_000000000000", -- twrite, gr3
  37 => b"00010_0010_01_000000000000", -- add, gr2
  38 => b"00000_0000_00_000000000001", -- 1
  39 => b"10000_0010_00_000000000000", -- tpoint, gr2
  40 => b"01111_0000_00_000000000000", -- tread, gr0
  41 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  42 => b"00111_0000_01_000000000000", -- bne
  43 => b"00000_0000_00_000000110101", -- E1LEFT
  44 => b"01110_0011_00_000000000000", -- twrite, gr3
  45 => b"00010_0010_01_000000000000", -- add, gr2
  46 => b"00000_0000_00_000000000001", -- 1
  47 => b"10000_0010_00_000000000000", -- tpoint, gr2
  48 => b"01111_0000_00_000000000000", -- tread, gr0
  49 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  50 => b"00111_0000_01_000000000000", -- bne
  51 => b"00000_0000_00_000000110101", -- E1LEFT
  52 => b"01110_0011_00_000000000000", -- twrite, gr3
  53 => b"00000_0010_00_001010101010", -- load, gr2, P1EXPLOSION1POS
  54 => b"00011_0010_01_000000000000", -- sub, gr2
  55 => b"00000_0000_00_000000000001", -- 1
  56 => b"10000_0010_00_000000000000", -- tpoint, gr2
  57 => b"01111_0000_00_000000000000", -- tread, gr0
  58 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  59 => b"00111_0000_01_000000000000", -- bne
  60 => b"00000_0000_00_000001000110", -- E1DOWN
  61 => b"01110_0011_00_000000000000", -- twrite, gr3
  62 => b"00011_0010_01_000000000000", -- sub, gr2
  63 => b"00000_0000_00_000000000001", -- 1
  64 => b"10000_0010_00_000000000000", -- tpoint, gr2
  65 => b"01111_0000_00_000000000000", -- tread, gr0
  66 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  67 => b"00111_0000_01_000000000000", -- bne
  68 => b"00000_0000_00_000001000110", -- E1DOWN
  69 => b"01110_0011_00_000000000000", -- twrite, gr3
  70 => b"00000_0010_00_001010101010", -- load, gr2, P1EXPLOSION1POS
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000001111", -- 15
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0000_00_000000000000", -- tread, gr0
  75 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  76 => b"00111_0000_01_000000000000", -- bne
  77 => b"00000_0000_00_000001010111", -- E1UP
  78 => b"01110_0011_00_000000000000", -- twrite, gr3
  79 => b"00010_0010_01_000000000000", -- add, gr2
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"10000_0010_00_000000000000", -- tpoint, gr2
  82 => b"01111_0000_00_000000000000", -- tread, gr0
  83 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  84 => b"00111_0000_01_000000000000", -- bne
  85 => b"00000_0000_00_000001010111", -- E1UP
  86 => b"01110_0011_00_000000000000", -- twrite, gr3
  87 => b"00000_0010_00_001010101010", -- load, gr2, P1EXPLOSION1POS
  88 => b"00011_0010_01_000000000000", -- sub, gr2
  89 => b"00000_0000_00_000000001111", -- 15
  90 => b"10000_0010_00_000000000000", -- tpoint, gr2
  91 => b"01111_0000_00_000000000000", -- tread, gr0
  92 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
  93 => b"00111_0000_01_000000000000", -- bne
  94 => b"00000_0000_00_000000001100", -- BOOM1_R
  95 => b"01110_0011_00_000000000000", -- twrite, gr3
  96 => b"00011_0010_01_000000000000", -- sub, gr2
  97 => b"00000_0000_00_000000001111", -- 15
  98 => b"10000_0010_00_000000000000", -- tpoint, gr2
  99 => b"01111_0000_00_000000000000", -- tread, gr0
 100 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 101 => b"00111_0000_01_000000000000", -- bne
 102 => b"00000_0000_00_000000001100", -- BOOM1_R
 103 => b"01110_0011_00_000000000000", -- twrite, gr3
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000000001100", -- BOOM1_R
 106 => b"00000_0000_00_001010111011", -- load, gr0, P2EXPLOSION1ACTIVE
 107 => b"00011_0000_01_000000000000", -- sub, gr0
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00111_0000_01_000000000000", -- bne
 110 => b"00000_0000_00_000000001110", -- BOOM2_R
 111 => b"00000_0000_00_001010111010", -- load, gr0, P2EXPLOSION1TIME
 112 => b"00011_0000_01_000000000000", -- sub, gr0
 113 => b"00000_0000_00_000000000001", -- 1
 114 => b"00001_0000_10_001010111010", -- store, gr0, P2EXPLOSION1TIME
 115 => b"00000_0000_00_001010111010", -- load, gr0, P2EXPLOSION1TIME
 116 => b"00011_0000_01_000000000000", -- sub, gr0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00111_0000_01_000000000000", -- bne
 119 => b"00000_0000_00_000000001110", -- BOOM2_R
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001010111011", -- store, gr0, P2EXPLOSION1ACTIVE
 123 => b"00000_0010_00_001010111100", -- load, gr2, P2EXPLOSION1POS
 124 => b"00000_0011_00_001011010011", -- load, gr3, GRASS
 125 => b"10000_0010_00_000000000000", -- tpoint, gr2
 126 => b"01110_0011_00_000000000000", -- twrite, gr3
 127 => b"00010_0010_01_000000000000", -- add, gr2
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"10000_0010_00_000000000000", -- tpoint, gr2
 130 => b"01111_0000_00_000000000000", -- tread, gr0
 131 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 132 => b"00111_0000_01_000000000000", -- bne
 133 => b"00000_0000_00_000010001111", -- E2LEFT
 134 => b"01110_0011_00_000000000000", -- twrite, gr3
 135 => b"00010_0010_01_000000000000", -- add, gr2
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0010_00_000000000000", -- tpoint, gr2
 138 => b"01111_0000_00_000000000000", -- tread, gr0
 139 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000010001111", -- E2LEFT
 142 => b"01110_0011_00_000000000000", -- twrite, gr3
 143 => b"00000_0010_00_001010111100", -- load, gr2, P2EXPLOSION1POS
 144 => b"00011_0010_01_000000000000", -- sub, gr2
 145 => b"00000_0000_00_000000000001", -- 1
 146 => b"10000_0010_00_000000000000", -- tpoint, gr2
 147 => b"01111_0000_00_000000000000", -- tread, gr0
 148 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 149 => b"00111_0000_01_000000000000", -- bne
 150 => b"00000_0000_00_000010100000", -- E2DOWN
 151 => b"01110_0011_00_000000000000", -- twrite, gr3
 152 => b"00011_0010_01_000000000000", -- sub, gr2
 153 => b"00000_0000_00_000000000001", -- 1
 154 => b"10000_0010_00_000000000000", -- tpoint, gr2
 155 => b"01111_0000_00_000000000000", -- tread, gr0
 156 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000010100000", -- E2DOWN
 159 => b"01110_0011_00_000000000000", -- twrite, gr3
 160 => b"00000_0010_00_001010111100", -- load, gr2, P2EXPLOSION1POS
 161 => b"00010_0010_01_000000000000", -- add, gr2
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"10000_0010_00_000000000000", -- tpoint, gr2
 164 => b"01111_0000_00_000000000000", -- tread, gr0
 165 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 166 => b"00111_0000_01_000000000000", -- bne
 167 => b"00000_0000_00_000010110001", -- E2UP
 168 => b"01110_0011_00_000000000000", -- twrite, gr3
 169 => b"00010_0010_01_000000000000", -- add, gr2
 170 => b"00000_0000_00_000000001111", -- 15
 171 => b"10000_0010_00_000000000000", -- tpoint, gr2
 172 => b"01111_0000_00_000000000000", -- tread, gr0
 173 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000010110001", -- E2UP
 176 => b"01110_0011_00_000000000000", -- twrite, gr3
 177 => b"00000_0010_00_001010111100", -- load, gr2, P2EXPLOSION1POS
 178 => b"00011_0010_01_000000000000", -- sub, gr2
 179 => b"00000_0000_00_000000001111", -- 15
 180 => b"10000_0010_00_000000000000", -- tpoint, gr2
 181 => b"01111_0000_00_000000000000", -- tread, gr0
 182 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 183 => b"00111_0000_01_000000000000", -- bne
 184 => b"00000_0000_00_000000001110", -- BOOM2_R
 185 => b"01110_0011_00_000000000000", -- twrite, gr3
 186 => b"00011_0010_01_000000000000", -- sub, gr2
 187 => b"00000_0000_00_000000001111", -- 15
 188 => b"10000_0010_00_000000000000", -- tpoint, gr2
 189 => b"01111_0000_00_000000000000", -- tread, gr0
 190 => b"00011_0000_00_001011010110", -- sub, gr0, EXPLOSION
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000001110", -- BOOM2_R
 193 => b"01110_0011_00_000000000000", -- twrite, gr3
 194 => b"00100_0000_01_000000000000", -- jump
 195 => b"00000_0000_00_000000001110", -- BOOM2_R
 196 => b"00000_0000_00_001010100111", -- load, gr0, P1BOMB1ACTIVE
 197 => b"00011_0000_01_000000000000", -- sub, gr0
 198 => b"00000_0000_00_000000000001", -- 1
 199 => b"00111_0000_01_000000000000", -- bne
 200 => b"00000_0000_00_000011010010", -- P2BOMB1
 201 => b"00000_0000_00_001010100110", -- load, gr0, P1BOMB1TIME
 202 => b"00011_0000_01_000000000000", -- sub, gr0
 203 => b"00000_0000_00_000000000001", -- 1
 204 => b"00001_0000_10_001010100110", -- store, gr0, P1BOMB1TIME
 205 => b"00000_0000_01_000000000000", -- load, gr0
 206 => b"00000_0000_00_000000000000", -- 0
 207 => b"00011_0000_00_001010100110", -- sub, gr0, P1BOMB1TIME
 208 => b"00110_0000_01_000000000000", -- beq
 209 => b"00000_0000_00_000011100010", -- P1EXPLOSION1INIT
 210 => b"00000_0000_00_001010111001", -- load, gr0, P2BOMB1ACTIVE
 211 => b"00011_0000_01_000000000000", -- sub, gr0
 212 => b"00000_0000_00_000000000001", -- 1
 213 => b"00111_0000_01_000000000000", -- bne
 214 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 215 => b"00000_0000_00_001010111000", -- load, gr0, P2BOMB1TIME
 216 => b"00011_0000_01_000000000000", -- sub, gr0
 217 => b"00000_0000_00_000000000001", -- 1
 218 => b"00001_0000_10_001010111000", -- store, gr0, P2BOMB1TIME
 219 => b"00000_0000_01_000000000000", -- load, gr0
 220 => b"00000_0000_00_000000000000", -- 0
 221 => b"00011_0000_00_001010111000", -- sub, gr0, P2BOMB1TIME
 222 => b"00110_0000_01_000000000000", -- beq
 223 => b"00000_0000_00_000011110001", -- P2EXPLOSION1INIT
 224 => b"00100_0000_01_000000000000", -- jump
 225 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 226 => b"00000_0000_00_001010100101", -- load, gr0, P1BOMB1POS
 227 => b"00001_0000_10_001010101010", -- store, gr0, P1EXPLOSION1POS
 228 => b"00000_0000_01_000000000000", -- load, gr0
 229 => b"00000_0000_00_000000000001", -- 1
 230 => b"00001_0000_10_001010101001", -- store, gr0, P1EXPLOSION1ACTIVE
 231 => b"00000_0000_01_000000000000", -- load, gr0
 232 => b"00000_0000_00_000000000010", -- 2
 233 => b"00001_0000_10_001010101000", -- store, gr0, P1EXPLOSION1TIME
 234 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 235 => b"00011_0000_01_000000000000", -- sub, gr0
 236 => b"00000_0000_00_000000000001", -- 1
 237 => b"00001_0000_10_001011001001", -- store, gr0, P1BOMBCOUNT
 238 => b"00000_0100_00_001010100101", -- load, gr4, P1BOMB1POS
 239 => b"00100_0000_01_000000000000", -- jump
 240 => b"00000_0000_00_000100000000", -- EXPLODE
 241 => b"00000_0000_00_001010110111", -- load, gr0, P2BOMB1POS
 242 => b"00001_0000_10_001010111100", -- store, gr0, P2EXPLOSION1POS
 243 => b"00000_0000_01_000000000000", -- load, gr0
 244 => b"00000_0000_00_000000000001", -- 1
 245 => b"00001_0000_10_001010111011", -- store, gr0, P2EXPLOSION1ACTIVE
 246 => b"00000_0000_01_000000000000", -- load, gr0
 247 => b"00000_0000_00_000000000010", -- 2
 248 => b"00001_0000_10_001010111010", -- store, gr0, P2EXPLOSION1TIME
 249 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 250 => b"00011_0000_01_000000000000", -- sub, gr0
 251 => b"00000_0000_00_000000000001", -- 1
 252 => b"00001_0000_10_001011001010", -- store, gr0, P2BOMBCOUNT
 253 => b"00000_0100_00_001010110111", -- load, gr4, P2BOMB1POS
 254 => b"00100_0000_01_000000000000", -- jump
 255 => b"00000_0000_00_000100000000", -- EXPLODE
 256 => b"00001_0100_10_001011010000", -- store, gr4, MOVE
 257 => b"00000_0010_00_001011010000", -- load, gr2, MOVE
 258 => b"00000_0011_00_001011010110", -- load, gr3, EXPLOSION
 259 => b"10000_0010_00_000000000000", -- tpoint, gr2
 260 => b"01110_0011_00_000000000000", -- twrite, gr3
 261 => b"00010_0010_01_000000000000", -- add, gr2
 262 => b"00000_0000_00_000000000001", -- 1
 263 => b"10000_0010_00_000000000000", -- tpoint, gr2
 264 => b"01111_0000_00_000000000000", -- tread, gr0
 265 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 266 => b"00110_0000_01_000000000000", -- beq
 267 => b"00000_0000_00_000100010101", -- EXPLODELEFT
 268 => b"01110_0011_00_000000000000", -- twrite, gr3
 269 => b"00010_0010_01_000000000000", -- add, gr2
 270 => b"00000_0000_00_000000000001", -- 1
 271 => b"10000_0010_00_000000000000", -- tpoint, gr2
 272 => b"01111_0000_00_000000000000", -- tread, gr0
 273 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 274 => b"00110_0000_01_000000000000", -- beq
 275 => b"00000_0000_00_000100010101", -- EXPLODELEFT
 276 => b"01110_0011_00_000000000000", -- twrite, gr3
 277 => b"00001_0100_10_001011010000", -- store, gr4, MOVE
 278 => b"00000_0010_00_001011010000", -- load, gr2, MOVE
 279 => b"00011_0010_01_000000000000", -- sub, gr2
 280 => b"00000_0000_00_000000000001", -- 1
 281 => b"10000_0010_00_000000000000", -- tpoint, gr2
 282 => b"01111_0000_00_000000000000", -- tread, gr0
 283 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 284 => b"00110_0000_01_000000000000", -- beq
 285 => b"00000_0000_00_000100100111", -- EXPLODEDOWN
 286 => b"01110_0011_00_000000000000", -- twrite, gr3
 287 => b"00011_0010_01_000000000000", -- sub, gr2
 288 => b"00000_0000_00_000000000001", -- 1
 289 => b"10000_0010_00_000000000000", -- tpoint, gr2
 290 => b"01111_0000_00_000000000000", -- tread, gr0
 291 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 292 => b"00110_0000_01_000000000000", -- beq
 293 => b"00000_0000_00_000100100111", -- EXPLODEDOWN
 294 => b"01110_0011_00_000000000000", -- twrite, gr3
 295 => b"00001_0100_10_001011010000", -- store, gr4, MOVE
 296 => b"00000_0010_00_001011010000", -- load, gr2, MOVE
 297 => b"00010_0010_01_000000000000", -- add, gr2
 298 => b"00000_0000_00_000000001111", -- 15
 299 => b"10000_0010_00_000000000000", -- tpoint, gr2
 300 => b"01111_0000_00_000000000000", -- tread, gr0
 301 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 302 => b"00110_0000_01_000000000000", -- beq
 303 => b"00000_0000_00_000100111001", -- EXPLODEUP
 304 => b"01110_0011_00_000000000000", -- twrite, gr3
 305 => b"00010_0010_01_000000000000", -- add, gr2
 306 => b"00000_0000_00_000000001111", -- 15
 307 => b"10000_0010_00_000000000000", -- tpoint, gr2
 308 => b"01111_0000_00_000000000000", -- tread, gr0
 309 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 310 => b"00110_0000_01_000000000000", -- beq
 311 => b"00000_0000_00_000100111001", -- EXPLODEUP
 312 => b"01110_0011_00_000000000000", -- twrite, gr3
 313 => b"00001_0100_10_001011010000", -- store, gr4, MOVE
 314 => b"00000_0010_00_001011010000", -- load, gr2, MOVE
 315 => b"00011_0010_01_000000000000", -- sub, gr2
 316 => b"00000_0000_00_000000001111", -- 15
 317 => b"10000_0010_00_000000000000", -- tpoint, gr2
 318 => b"01111_0000_00_000000000000", -- tread, gr0
 319 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 320 => b"00110_0000_01_000000000000", -- beq
 321 => b"00000_0000_00_000011000100", -- TICKBOMBS
 322 => b"01110_0011_00_000000000000", -- twrite, gr3
 323 => b"00011_0010_01_000000000000", -- sub, gr2
 324 => b"00000_0000_00_000000001111", -- 15
 325 => b"10000_0010_00_000000000000", -- tpoint, gr2
 326 => b"01111_0000_00_000000000000", -- tread, gr0
 327 => b"00011_0000_00_001011010100", -- sub, gr0, WALL
 328 => b"00110_0000_01_000000000000", -- beq
 329 => b"00000_0000_00_000011000100", -- TICKBOMBS
 330 => b"01110_0011_00_000000000000", -- twrite, gr3
 331 => b"00100_0000_01_000000000000", -- jump
 332 => b"00000_0000_00_000011000100", -- TICKBOMBS
 333 => b"10101_0000_01_000000000000", -- btn1
 334 => b"00000_0000_00_000101010011", -- BTN1
 335 => b"11010_0000_01_000000000000", -- btn2
 336 => b"00000_0000_00_000110101101", -- BTN2
 337 => b"00100_0000_01_000000000000", -- jump
 338 => b"00000_0000_00_000000000100", -- BUTTON_R
 339 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 340 => b"00011_0000_00_001011001011", -- sub, gr0, MAXBOMBS
 341 => b"00110_0000_01_000000000000", -- beq
 342 => b"00000_0000_00_000101001111", -- BTN1_R
 343 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 344 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 345 => b"00000_0000_00_001011001101", -- load, gr0, YPOS1
 346 => b"01000_0000_01_000000000000", -- mul, gr0
 347 => b"00000_0000_00_000000001111", -- 15
 348 => b"00010_0000_00_001011001100", -- add, gr0, XPOS1
 349 => b"10000_0000_00_000000000000", -- tpoint, gr0
 350 => b"01111_0001_00_000000000000", -- tread, gr1
 351 => b"00011_0001_00_001011010111", -- sub, gr1, EGG
 352 => b"00110_0000_01_000000000000", -- beq
 353 => b"00000_0000_00_000101001111", -- BTN1_R
 354 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 355 => b"00011_0000_01_000000000000", -- sub, gr0
 356 => b"00000_0000_00_000000000000", -- 0
 357 => b"00110_0000_01_000000000000", -- beq
 358 => b"00000_0000_00_000101110111", -- P1PLACEBOMB1
 359 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 360 => b"00011_0000_01_000000000000", -- sub, gr0
 361 => b"00000_0000_00_000000000001", -- 1
 362 => b"00110_0000_01_000000000000", -- beq
 363 => b"00000_0000_00_000110001001", -- P1PLACEBOMB2
 364 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 365 => b"00011_0000_01_000000000000", -- sub, gr0
 366 => b"00000_0000_00_000000000010", -- 2
 367 => b"00110_0000_01_000000000000", -- beq
 368 => b"00000_0000_00_000110001001", -- P1PLACEBOMB2
 369 => b"00000_0000_00_001011001001", -- load, gr0, P1BOMBCOUNT
 370 => b"00010_0000_01_000000000000", -- add, gr0
 371 => b"00000_0000_00_000000000001", -- 1
 372 => b"00001_0000_10_001011001001", -- store, gr0, P1BOMBCOUNT
 373 => b"00100_0000_01_000000000000", -- jump
 374 => b"00000_0000_00_000101001111", -- BTN1_R
 375 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 376 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 377 => b"00000_0011_00_001011001101", -- load, gr3, YPOS1
 378 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 379 => b"01000_0011_01_000000000000", -- mul, gr3
 380 => b"00000_0000_00_000000001111", -- 15
 381 => b"00010_0011_00_001011001100", -- add, gr3, XPOS1
 382 => b"10000_0011_00_000000000000", -- tpoint, gr3
 383 => b"01110_0010_00_000000000000", -- twrite, gr2
 384 => b"00000_0000_01_000000000000", -- load, gr0
 385 => b"00000_0000_00_000000000001", -- 1
 386 => b"00001_0000_10_001010100111", -- store, gr0, P1BOMB1ACTIVE
 387 => b"00001_0011_10_001010100101", -- store, gr3, P1BOMB1POS
 388 => b"00000_0000_01_000000000000", -- load, gr0
 389 => b"00000_0000_00_000000010000", -- 16
 390 => b"00001_0000_10_001010100110", -- store, gr0, P1BOMB1TIME
 391 => b"00100_0000_01_000000000000", -- jump
 392 => b"00000_0000_00_000101110001", -- P1INCREASEBOMBCOUNTER
 393 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 394 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 395 => b"00000_0011_00_001011001101", -- load, gr3, YPOS1
 396 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 397 => b"01000_0011_01_000000000000", -- mul, gr3
 398 => b"00000_0000_00_000000001111", -- 15
 399 => b"00010_0011_00_001011001100", -- add, gr3, XPOS1
 400 => b"10000_0011_00_000000000000", -- tpoint, gr3
 401 => b"01110_0010_00_000000000000", -- twrite, gr2
 402 => b"00000_0000_01_000000000000", -- load, gr0
 403 => b"00000_0000_00_000000000001", -- 1
 404 => b"00001_0000_10_001010101101", -- store, gr0, P1BOMB2ACTIVE
 405 => b"00001_0011_10_001010101011", -- store, gr3, P1BOMB2POS
 406 => b"00000_0000_01_000000000000", -- load, gr0
 407 => b"00000_0000_00_000000010000", -- 16
 408 => b"00001_0000_10_001010101100", -- store, gr0, P1BOMB2TIME
 409 => b"00100_0000_01_000000000000", -- jump
 410 => b"00000_0000_00_000101110001", -- P1INCREASEBOMBCOUNTER
 411 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 412 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 413 => b"00000_0011_00_001011001101", -- load, gr3, YPOS1
 414 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 415 => b"01000_0011_01_000000000000", -- mul, gr3
 416 => b"00000_0000_00_000000001111", -- 15
 417 => b"00010_0011_00_001011001100", -- add, gr3, XPOS1
 418 => b"10000_0011_00_000000000000", -- tpoint, gr3
 419 => b"01110_0010_00_000000000000", -- twrite, gr2
 420 => b"00000_0000_01_000000000000", -- load, gr0
 421 => b"00000_0000_00_000000000001", -- 1
 422 => b"00001_0000_10_001010110011", -- store, gr0, P1BOMB3ACTIVE
 423 => b"00001_0011_10_001010110001", -- store, gr3, P1BOMB3POS
 424 => b"00000_0000_01_000000000000", -- load, gr0
 425 => b"00000_0000_00_000000010000", -- 16
 426 => b"00001_0000_10_001010110010", -- store, gr0, P1BOMB3TIME
 427 => b"00100_0000_01_000000000000", -- jump
 428 => b"00000_0000_00_000101110001", -- P1INCREASEBOMBCOUNTER
 429 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 430 => b"00011_0000_00_001011001011", -- sub, gr0, MAXBOMBS
 431 => b"00110_0000_01_000000000000", -- beq
 432 => b"00000_0000_00_000101010001", -- BTN2_R
 433 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 434 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 435 => b"00000_0000_00_001011001111", -- load, gr0, YPOS2
 436 => b"01000_0000_01_000000000000", -- mul, gr0
 437 => b"00000_0000_00_000000001111", -- 15
 438 => b"00010_0000_00_001011001110", -- add, gr0, XPOS2
 439 => b"10000_0000_00_000000000000", -- tpoint, gr0
 440 => b"01111_0001_00_000000000000", -- tread, gr1
 441 => b"00011_0001_00_001011010111", -- sub, gr1, EGG
 442 => b"00110_0000_01_000000000000", -- beq
 443 => b"00000_0000_00_000101010001", -- BTN2_R
 444 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 445 => b"00011_0000_01_000000000000", -- sub, gr0
 446 => b"00000_0000_00_000000000000", -- 0
 447 => b"00110_0000_01_000000000000", -- beq
 448 => b"00000_0000_00_000111010001", -- P2PLACEBOMB1
 449 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 450 => b"00011_0000_01_000000000000", -- sub, gr0
 451 => b"00000_0000_00_000000000001", -- 1
 452 => b"00110_0000_01_000000000000", -- beq
 453 => b"00000_0000_00_000111100011", -- P2PLACEBOMB2
 454 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 455 => b"00011_0000_01_000000000000", -- sub, gr0
 456 => b"00000_0000_00_000000000010", -- 2
 457 => b"00110_0000_01_000000000000", -- beq
 458 => b"00000_0000_00_000111110101", -- P2PLACEBOMB3
 459 => b"00000_0000_00_001011001010", -- load, gr0, P2BOMBCOUNT
 460 => b"00010_0000_01_000000000000", -- add, gr0
 461 => b"00000_0000_00_000000000001", -- 1
 462 => b"00001_0000_10_001011001010", -- store, gr0, P2BOMBCOUNT
 463 => b"00100_0000_01_000000000000", -- jump
 464 => b"00000_0000_00_000101010001", -- BTN2_R
 465 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 466 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 467 => b"00000_0011_00_001011001111", -- load, gr3, YPOS2
 468 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 469 => b"01000_0011_01_000000000000", -- mul, gr3
 470 => b"00000_0000_00_000000001111", -- 15
 471 => b"00010_0011_00_001011001110", -- add, gr3, XPOS2
 472 => b"10000_0011_00_000000000000", -- tpoint, gr3
 473 => b"01110_0010_00_000000000000", -- twrite, gr2
 474 => b"00000_0000_01_000000000000", -- load, gr0
 475 => b"00000_0000_00_000000000001", -- 1
 476 => b"00001_0000_10_001010111001", -- store, gr0, P2BOMB1ACTIVE
 477 => b"00001_0011_10_001010110111", -- store, gr3, P2BOMB1POS
 478 => b"00000_0000_01_000000000000", -- load, gr0
 479 => b"00000_0000_00_000000010000", -- 16
 480 => b"00001_0000_10_001010111000", -- store, gr0, P2BOMB1TIME
 481 => b"00100_0000_01_000000000000", -- jump
 482 => b"00000_0000_00_000111001011", -- P2INCREASEBOMBCOUNTER
 483 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 484 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 485 => b"00000_0011_00_001011001111", -- load, gr3, YPOS2
 486 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 487 => b"01000_0011_01_000000000000", -- mul, gr3
 488 => b"00000_0000_00_000000001111", -- 15
 489 => b"00010_0011_00_001011001110", -- add, gr3, XPOS2
 490 => b"10000_0011_00_000000000000", -- tpoint, gr3
 491 => b"01110_0010_00_000000000000", -- twrite, gr2
 492 => b"00000_0000_01_000000000000", -- load, gr0
 493 => b"00000_0000_00_000000000001", -- 1
 494 => b"00001_0000_10_001010111111", -- store, gr0, P2BOMB2ACTIVE
 495 => b"00001_0011_10_001010111101", -- store, gr3, P2BOMB2POS
 496 => b"00000_0000_01_000000000000", -- load, gr0
 497 => b"00000_0000_00_000000010000", -- 16
 498 => b"00001_0000_10_001010111110", -- store, gr0, P2BOMB2TIME
 499 => b"00100_0000_01_000000000000", -- jump
 500 => b"00000_0000_00_000111001011", -- P2INCREASEBOMBCOUNTER
 501 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 502 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 503 => b"00000_0011_00_001011001111", -- load, gr3, YPOS2
 504 => b"00000_0010_00_001011010111", -- load, gr2, EGG
 505 => b"01000_0011_01_000000000000", -- mul, gr3
 506 => b"00000_0000_00_000000001111", -- 15
 507 => b"00010_0011_00_001011001110", -- add, gr3, XPOS2
 508 => b"10000_0011_00_000000000000", -- tpoint, gr3
 509 => b"01110_0010_00_000000000000", -- twrite, gr2
 510 => b"00000_0000_01_000000000000", -- load, gr0
 511 => b"00000_0000_00_000000000001", -- 1
 512 => b"00001_0000_10_001011000101", -- store, gr0, P2BOMB3ACTIVE
 513 => b"00001_0011_10_001011000011", -- store, gr3, P2BOMB3POS
 514 => b"00000_0000_01_000000000000", -- load, gr0
 515 => b"00000_0000_00_000000010000", -- 16
 516 => b"00001_0000_10_001011000100", -- store, gr0, P2BOMB3TIME
 517 => b"00100_0000_01_000000000000", -- jump
 518 => b"00000_0000_00_000111001011", -- P2INCREASEBOMBCOUNTER
 519 => b"00100_0000_01_000000000000", -- jump
 520 => b"00000_0000_00_001010100011", -- COUNT1
 521 => b"10001_0000_01_000000000000", -- joy1r
 522 => b"00000_0000_00_001000011011", -- P1R
 523 => b"10011_0000_01_000000000000", -- joy1l
 524 => b"00000_0000_00_001000111101", -- P1L
 525 => b"10010_0000_01_000000000000", -- joy1u
 526 => b"00000_0000_00_001000101100", -- P1U
 527 => b"10100_0000_01_000000000000", -- joy1d
 528 => b"00000_0000_00_001001001110", -- P1D
 529 => b"10110_0000_01_000000000000", -- joy2r
 530 => b"00000_0000_00_001001011111", -- P2R
 531 => b"11000_0000_01_000000000000", -- joy2l
 532 => b"00000_0000_00_001010000001", -- P2L
 533 => b"10111_0000_01_000000000000", -- joy2u
 534 => b"00000_0000_00_001001110000", -- P2U
 535 => b"11001_0000_01_000000000000", -- joy2d
 536 => b"00000_0000_00_001010010010", -- P2D
 537 => b"00100_0000_01_000000000000", -- jump
 538 => b"00000_0000_00_000000000010", -- CONTROL_R
 539 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 540 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 541 => b"00000_0000_00_001011001101", -- load, gr0, YPOS1
 542 => b"01000_0000_01_000000000000", -- mul, gr0
 543 => b"00000_0000_00_000000001111", -- 15
 544 => b"00010_0000_00_001011001100", -- add, gr0, XPOS1
 545 => b"00010_0000_01_000000000000", -- add, gr0
 546 => b"00000_0000_00_000000000001", -- 1
 547 => b"10000_0000_00_000000000000", -- tpoint, gr0
 548 => b"01111_0001_00_000000000000", -- tread, gr1
 549 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 550 => b"00111_0000_01_000000000000", -- bne
 551 => b"00000_0000_00_001000001101", -- J1
 552 => b"00010_1100_01_000000000000", -- add, gr12
 553 => b"00000_0000_00_000000000001", -- 1
 554 => b"00100_0000_01_000000000000", -- jump
 555 => b"00000_0000_00_001000001101", -- J1
 556 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 557 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 558 => b"00000_0000_00_001011001101", -- load, gr0, YPOS1
 559 => b"00011_0000_01_000000000000", -- sub, gr0
 560 => b"00000_0000_00_000000000001", -- 1
 561 => b"01000_0000_01_000000000000", -- mul, gr0
 562 => b"00000_0000_00_000000001111", -- 15
 563 => b"00010_0000_00_001011001100", -- add, gr0, XPOS1
 564 => b"10000_0000_00_000000000000", -- tpoint, gr0
 565 => b"01111_0001_00_000000000000", -- tread, gr1
 566 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 567 => b"00111_0000_01_000000000000", -- bne
 568 => b"00000_0000_00_001000010001", -- J2
 569 => b"00011_1101_01_000000000000", -- sub, gr13
 570 => b"00000_0000_00_000000000001", -- 1
 571 => b"00100_0000_01_000000000000", -- jump
 572 => b"00000_0000_00_001000010001", -- J2
 573 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 574 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 575 => b"00000_0000_00_001011001101", -- load, gr0, YPOS1
 576 => b"01000_0000_01_000000000000", -- mul, gr0
 577 => b"00000_0000_00_000000001111", -- 15
 578 => b"00010_0000_00_001011001100", -- add, gr0, XPOS1
 579 => b"00011_0000_01_000000000000", -- sub, gr0
 580 => b"00000_0000_00_000000000001", -- 1
 581 => b"10000_0000_00_000000000000", -- tpoint, gr0
 582 => b"01111_0001_00_000000000000", -- tread, gr1
 583 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 584 => b"00111_0000_01_000000000000", -- bne
 585 => b"00000_0000_00_001000001101", -- J1
 586 => b"00011_1100_01_000000000000", -- sub, gr12
 587 => b"00000_0000_00_000000000001", -- 1
 588 => b"00100_0000_01_000000000000", -- jump
 589 => b"00000_0000_00_001000001101", -- J1
 590 => b"00001_1100_10_001011001100", -- store, gr12, XPOS1
 591 => b"00001_1101_10_001011001101", -- store, gr13, YPOS1
 592 => b"00000_0000_00_001011001101", -- load, gr0, YPOS1
 593 => b"00010_0000_01_000000000000", -- add, gr0
 594 => b"00000_0000_00_000000000001", -- 1
 595 => b"01000_0000_01_000000000000", -- mul, gr0
 596 => b"00000_0000_00_000000001111", -- 15
 597 => b"00010_0000_00_001011001100", -- add, gr0, XPOS1
 598 => b"10000_0000_00_000000000000", -- tpoint, gr0
 599 => b"01111_0001_00_000000000000", -- tread, gr1
 600 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 601 => b"00111_0000_01_000000000000", -- bne
 602 => b"00000_0000_00_001000010001", -- J2
 603 => b"00010_1101_01_000000000000", -- add, gr13
 604 => b"00000_0000_00_000000000001", -- 1
 605 => b"00100_0000_01_000000000000", -- jump
 606 => b"00000_0000_00_001000010001", -- J2
 607 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 608 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 609 => b"00000_0000_00_001011001111", -- load, gr0, YPOS2
 610 => b"01000_0000_01_000000000000", -- mul, gr0
 611 => b"00000_0000_00_000000001111", -- 15
 612 => b"00010_0000_00_001011001110", -- add, gr0, XPOS2
 613 => b"00010_0000_01_000000000000", -- add, gr0
 614 => b"00000_0000_00_000000000001", -- 1
 615 => b"10000_0000_00_000000000000", -- tpoint, gr0
 616 => b"01111_0001_00_000000000000", -- tread, gr1
 617 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 618 => b"00111_0000_01_000000000000", -- bne
 619 => b"00000_0000_00_001000010101", -- J3
 620 => b"00010_1110_01_000000000000", -- add, gr14
 621 => b"00000_0000_00_000000000001", -- 1
 622 => b"00100_0000_01_000000000000", -- jump
 623 => b"00000_0000_00_001000010101", -- J3
 624 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 625 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 626 => b"00000_0000_00_001011001111", -- load, gr0, YPOS2
 627 => b"00011_0000_01_000000000000", -- sub, gr0
 628 => b"00000_0000_00_000000000001", -- 1
 629 => b"01000_0000_01_000000000000", -- mul, gr0
 630 => b"00000_0000_00_000000001111", -- 15
 631 => b"00010_0000_00_001011001110", -- add, gr0, XPOS2
 632 => b"10000_0000_00_000000000000", -- tpoint, gr0
 633 => b"01111_0001_00_000000000000", -- tread, gr1
 634 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 635 => b"00111_0000_01_000000000000", -- bne
 636 => b"00000_0000_00_000000000010", -- CONTROL_R
 637 => b"00011_1111_01_000000000000", -- sub, gr15
 638 => b"00000_0000_00_000000000001", -- 1
 639 => b"00100_0000_01_000000000000", -- jump
 640 => b"00000_0000_00_000000000010", -- CONTROL_R
 641 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 642 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 643 => b"00000_0000_00_001011001111", -- load, gr0, YPOS2
 644 => b"01000_0000_01_000000000000", -- mul, gr0
 645 => b"00000_0000_00_000000001111", -- 15
 646 => b"00010_0000_00_001011001110", -- add, gr0, XPOS2
 647 => b"00011_0000_01_000000000000", -- sub, gr0
 648 => b"00000_0000_00_000000000001", -- 1
 649 => b"10000_0000_00_000000000000", -- tpoint, gr0
 650 => b"01111_0001_00_000000000000", -- tread, gr1
 651 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 652 => b"00111_0000_01_000000000000", -- bne
 653 => b"00000_0000_00_001000010101", -- J3
 654 => b"00011_1110_01_000000000000", -- sub, gr14
 655 => b"00000_0000_00_000000000001", -- 1
 656 => b"00100_0000_01_000000000000", -- jump
 657 => b"00000_0000_00_001000010101", -- J3
 658 => b"00001_1110_10_001011001110", -- store, gr14, XPOS2
 659 => b"00001_1111_10_001011001111", -- store, gr15, YPOS2
 660 => b"00000_0000_00_001011001111", -- load, gr0, YPOS2
 661 => b"00010_0000_01_000000000000", -- add, gr0
 662 => b"00000_0000_00_000000000001", -- 1
 663 => b"01000_0000_01_000000000000", -- mul, gr0
 664 => b"00000_0000_00_000000001111", -- 15
 665 => b"00010_0000_00_001011001110", -- add, gr0, XPOS2
 666 => b"10000_0000_00_000000000000", -- tpoint, gr0
 667 => b"01111_0001_00_000000000000", -- tread, gr1
 668 => b"00011_0001_00_001011010011", -- sub, gr1, GRASS
 669 => b"00111_0000_01_000000000000", -- bne
 670 => b"00000_0000_00_000000000010", -- CONTROL_R
 671 => b"00010_1111_01_000000000000", -- add, gr15
 672 => b"00000_0000_00_000000000001", -- 1
 673 => b"00100_0000_01_000000000000", -- jump
 674 => b"00000_0000_00_000000000010", -- CONTROL_R
 675 => b"00100_0000_01_000000000000", -- jump
 676 => b"00000_0000_00_001000001001", -- COUNT_R
 677 => b"00000_0000_00_000000000000", -- 0
 678 => b"00000_0000_00_000000000000", -- 0
 679 => b"00000_0000_00_000000000000", -- 0
 680 => b"00000_0000_00_000000000000", -- 0
 681 => b"00000_0000_00_000000000000", -- 0
 682 => b"00000_0000_00_000000000000", -- 0
 683 => b"00000_0000_00_000000000000", -- 0
 684 => b"00000_0000_00_000000000000", -- 0
 685 => b"00000_0000_00_000000000000", -- 0
 686 => b"00000_0000_00_000000000000", -- 0
 687 => b"00000_0000_00_000000000000", -- 0
 688 => b"00000_0000_00_000000000000", -- 0
 689 => b"00000_0000_00_000000000000", -- 0
 690 => b"00000_0000_00_000000000000", -- 0
 691 => b"00000_0000_00_000000000000", -- 0
 692 => b"00000_0000_00_000000000000", -- 0
 693 => b"00000_0000_00_000000000000", -- 0
 694 => b"00000_0000_00_000000000000", -- 0
 695 => b"00000_0000_00_000000000000", -- 0
 696 => b"00000_0000_00_000000000000", -- 0
 697 => b"00000_0000_00_000000000000", -- 0
 698 => b"00000_0000_00_000000000000", -- 0
 699 => b"00000_0000_00_000000000000", -- 0
 700 => b"00000_0000_00_000000000000", -- 0
 701 => b"00000_0000_00_000000000000", -- 0
 702 => b"00000_0000_00_000000000000", -- 0
 703 => b"00000_0000_00_000000000000", -- 0
 704 => b"00000_0000_00_000000000000", -- 0
 705 => b"00000_0000_00_000000000000", -- 0
 706 => b"00000_0000_00_000000000000", -- 0
 707 => b"00000_0000_00_000000000000", -- 0
 708 => b"00000_0000_00_000000000000", -- 0
 709 => b"00000_0000_00_000000000000", -- 0
 710 => b"00000_0000_00_000000000000", -- 0
 711 => b"00000_0000_00_000000000000", -- 0
 712 => b"00000_0000_00_000000000000", -- 0
 713 => b"00000_0000_00_000000000000", -- 0
 714 => b"00000_0000_00_000000000000", -- 0
 715 => b"00000_0000_00_000000000011", -- 3
 716 => b"00000_0000_00_000000000000", -- 0
 717 => b"00000_0000_00_000000000000", -- 0
 718 => b"00000_0000_00_000000000000", -- 0
 719 => b"00000_0000_00_000000000000", -- 0
 720 => b"00000_0000_00_000000000000", -- 0
 721 => b"00000_0000_00_000000000000", -- 0
 722 => b"00000_0000_00_000000000000", -- 0
 723 => b"00000_0000_00_000000000000", -- 0
 724 => b"00000_0000_00_000000000001", -- 1
 725 => b"00000_0000_00_000000000010", -- 2
 726 => b"00000_0000_00_000000000011", -- 3
 727 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
