library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00101_0000_01_000000000000", -- sleep
   1 => b"00000_0000_00_000000000001", -- 1
   2 => b"00000_0001_01_000000000000", -- load, gr1
   3 => b"00000_0000_00_000000010010", -- 18
   4 => b"00000_0010_01_000000000000", -- load, gr2
   5 => b"00000_0000_00_000000000100", -- 4
   6 => b"10000_0001_00_000000000000", -- tpoint, gr1
   7 => b"01110_0010_00_000000000000", -- twrite, gr2
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000101110", -- CONTROL
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000001110", -- BUTTON
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000000001000", -- MAIN
  14 => b"10101_0000_01_000000000000", -- btn1
  15 => b"00000_0000_00_000000010101", -- BTN1
  16 => b"11010_0000_01_000000000000", -- btn2
  17 => b"00000_0000_00_000000100001", -- BTN2
  18 => b"00100_0000_01_000000000000", -- jump
  19 => b"00000_0000_00_000000001100", -- BUTTON_R
  20 => b"00001_1100_10_000001110100", -- store, gr12, XPOS1
  21 => b"00001_1101_10_000001110101", -- store, gr13, YPOS1
  22 => b"00000_0011_00_000001110101", -- load, gr3, YPOS1
  23 => b"00000_0010_00_000001110011", -- load, gr2, EGG
  24 => b"00000_0000_00_000001110100", -- load, gr0, XPOS1
  25 => b"01000_0011_01_000000000000", -- mul, gr3
  26 => b"00000_0000_00_000000001111", -- 15
  27 => b"11011_0011_00_000000000000", -- addgr, gr3
  28 => b"00000_0000_00_000000000000", -- gr0
  29 => b"10000_0011_00_000000000000", -- tpoint, gr3
  30 => b"01110_0010_00_000000000000", -- twrite, gr2
  31 => b"00100_0000_01_000000000000", -- jump
  32 => b"00000_0000_00_000000010000", -- BTN1_R
  33 => b"00001_1110_10_000001110110", -- store, gr14, XPOS2
  34 => b"00001_1111_10_000001110111", -- store, gr15, YPOS2
  35 => b"00000_0011_00_000001110111", -- load, gr3, YPOS2
  36 => b"00000_0010_00_000001110011", -- load, gr2, EGG
  37 => b"00000_0000_00_000001110110", -- load, gr0, XPOS2
  38 => b"01000_0011_01_000000000000", -- mul, gr3
  39 => b"00000_0000_00_000000001111", -- 15
  40 => b"11011_0011_00_000000000000", -- addgr, gr3
  41 => b"10000_0011_00_000000000000", -- tpoint, gr3
  42 => b"01110_0010_00_000000000000", -- twrite, gr2
  43 => b"00100_0000_01_000000000000", -- jump
  44 => b"00000_0000_00_000000010010", -- BTN2_R
  45 => b"00000_0000_00_000000000000", -- 0
  46 => b"10001_0000_01_000000000000", -- joy1r
  47 => b"00000_0000_00_000000111111", -- P1R
  48 => b"10011_0000_01_000000000000", -- joy1l
  49 => b"00000_0000_00_000001010110", -- P1L
  50 => b"10010_0000_01_000000000000", -- joy1u
  51 => b"00000_0000_00_000001010010", -- P1U
  52 => b"10100_0000_01_000000000000", -- joy1d
  53 => b"00000_0000_00_000001011010", -- P1D
  54 => b"10110_0000_01_000000000000", -- joy2r
  55 => b"00000_0000_00_000001011110", -- P2R
  56 => b"11000_0000_01_000000000000", -- joy2l
  57 => b"00000_0000_00_000001100110", -- P2L
  58 => b"10111_0000_01_000000000000", -- joy2u
  59 => b"00000_0000_00_000001100010", -- P2U
  60 => b"11001_0000_01_000000000000", -- joy2d
  61 => b"00000_0000_00_000001101010", -- P2D
  62 => b"00100_0000_01_000000000000", -- jump
  63 => b"00000_0000_00_000000001010", -- CONTROL_R
  64 => b"00001_1101_10_000001110111", -- store, gr13, MOVE
  65 => b"00000_0010_00_000001110111", -- load, gr2, MOVE
  66 => b"00001_1100_10_000001110111", -- store, gr12, MOVE
  67 => b"00000_0000_00_000001110111", -- load, gr0, MOVE
  68 => b"01000_0010_01_000000000000", -- mul, gr2
  69 => b"00000_0000_00_000000001111", -- 15
  70 => b"11011_0010_00_000000000000", -- addgr, gr2
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000000001", -- 1
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0011_00_000000000000", -- tread, gr3
  75 => b"00011_0011_01_000000000000", -- sub, gr3
  76 => b"00000_0000_00_000000000000", -- 0
  77 => b"00111_0000_01_000000000000", -- bne
  78 => b"00000_0000_00_000000110001", -- J1
  79 => b"00010_1100_01_000000000000", -- add, gr12
  80 => b"00000_0000_00_000000000001", -- 1
  81 => b"00100_0000_01_000000000000", -- jump
  82 => b"00000_0000_00_000000110001", -- J1
  83 => b"00011_1101_01_000000000000", -- sub, gr13
  84 => b"00000_0000_00_000000000001", -- 1
  85 => b"00100_0000_01_000000000000", -- jump
  86 => b"00000_0000_00_000000110101", -- J2
  87 => b"00011_1100_01_000000000000", -- sub, gr12
  88 => b"00000_0000_00_000000000001", -- 1
  89 => b"00100_0000_01_000000000000", -- jump
  90 => b"00000_0000_00_000000110001", -- J1
  91 => b"00010_1101_01_000000000000", -- add, gr13
  92 => b"00000_0000_00_000000000001", -- 1
  93 => b"00100_0000_01_000000000000", -- jump
  94 => b"00000_0000_00_000000110101", -- J2
  95 => b"00010_1110_01_000000000000", -- add, gr14
  96 => b"00000_0000_00_000000000001", -- 1
  97 => b"00100_0000_01_000000000000", -- jump
  98 => b"00000_0000_00_000000111001", -- J3
  99 => b"00011_1111_01_000000000000", -- sub, gr15
 100 => b"00000_0000_00_000000000001", -- 1
 101 => b"00100_0000_01_000000000000", -- jump
 102 => b"00000_0000_00_000000001010", -- CONTROL_R
 103 => b"00011_1110_01_000000000000", -- sub, gr14
 104 => b"00000_0000_00_000000000001", -- 1
 105 => b"00100_0000_01_000000000000", -- jump
 106 => b"00000_0000_00_000000111001", -- J3
 107 => b"00010_1111_01_000000000000", -- add, gr15
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00100_0000_01_000000000000", -- jump
 110 => b"00000_0000_00_000000001010", -- CONTROL_R
 111 => b"00000_0000_00_000000000000", -- 0
 112 => b"00000_0000_00_000000000001", -- 1
 113 => b"00000_0000_00_000000000010", -- 2
 114 => b"00000_0000_00_000000000011", -- 3
 115 => b"00000_0000_00_000000000100", -- 4
 116 => b"00000_0000_00_000000000000", -- 0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00000_0000_00_000000000000", -- 0
 119 => b"00000_0000_00_000000000000", -- 0
 120 => b"00000_0000_00_000000000000", -- 0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00000_0000_00_000000000000", -- 0





    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


