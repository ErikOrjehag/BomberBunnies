library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_0000_01_000000000000", -- load, gr0
   1 => b"00000_0000_00_000000000000", -- 0
   2 => b"00001_0000_10_010000100110", -- store, gr0, P1DEAD
   3 => b"00001_0000_10_010000100111", -- store, gr0, P2DEAD
   4 => b"00001_0000_10_010001001100", -- store, gr0, P1BOMBCOUNT
   5 => b"00001_0000_10_010001001101", -- store, gr0, P2BOMBCOUNT
   6 => b"00000_1100_01_000000000000", -- load, gr12
   7 => b"00000_0000_00_000000000001", -- 1
   8 => b"00000_1101_01_000000000000", -- load, gr13
   9 => b"00000_0000_00_000000000001", -- 1
  10 => b"00000_1110_01_000000000000", -- load, gr14
  11 => b"00000_0000_00_000000001101", -- 13
  12 => b"00000_1111_01_000000000000", -- load, gr15
  13 => b"00000_0000_00_000000001011", -- 11
  14 => b"00001_0000_10_010000101000", -- store, gr0, P1BOMB1POS
  15 => b"00001_0000_10_010000101010", -- store, gr0, P1BOMB1ACTIVE
  16 => b"00001_0000_10_010000101001", -- store, gr0, P1BOMB1TIME
  17 => b"00001_0000_10_010000101110", -- store, gr0, P1BOMB2POS
  18 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMB2ACTIVE
  19 => b"00001_0000_10_010000101111", -- store, gr0, P1BOMB2TIME
  20 => b"00001_0000_10_010000110100", -- store, gr0, P1BOMB3POS
  21 => b"00001_0000_10_010000110110", -- store, gr0, P1BOMB3ACTIVE
  22 => b"00001_0000_10_010000110101", -- store, gr0, P1BOMB3TIME
  23 => b"00001_0000_10_010000111010", -- store, gr0, P2BOMB1POS
  24 => b"00001_0000_10_010000111100", -- store, gr0, P2BOMB1ACTIVE
  25 => b"00001_0000_10_010000111011", -- store, gr0, P2BOMB1TIME
  26 => b"00001_0000_10_010001000000", -- store, gr0, P2BOMB2POS
  27 => b"00001_0000_10_010001000010", -- store, gr0, P2BOMB2ACTIVE
  28 => b"00001_0000_10_010001000001", -- store, gr0, P2BOMB2TIME
  29 => b"00001_0000_10_010001000110", -- store, gr0, P2BOMB3POS
  30 => b"00001_0000_10_010001001000", -- store, gr0, P2BOMB3ACTIVE
  31 => b"00001_0000_10_010001000111", -- store, gr0, P2BOMB3TIME
  32 => b"00001_0000_10_010000101101", -- store, gr0, P1EXPLOSION1POS
  33 => b"00001_0000_10_010000101100", -- store, gr0, P1EXPLOSION1ACTIVE
  34 => b"00001_0000_10_010000101011", -- store, gr0, P1EXPLOSION1TIME
  35 => b"00001_0000_10_010000110011", -- store, gr0, P1EXPLOSION2POS
  36 => b"00001_0000_10_010000110010", -- store, gr0, P1EXPLOSION2ACTIVE
  37 => b"00001_0000_10_010000110001", -- store, gr0, P1EXPLOSION2TIME
  38 => b"00001_0000_10_010000111001", -- store, gr0, P1EXPLOSION3POS
  39 => b"00001_0000_10_010000111000", -- store, gr0, P1EXPLOSION3ACTIVE
  40 => b"00001_0000_10_010000110111", -- store, gr0, P1EXPLOSION3TIME
  41 => b"00001_0000_10_010000111111", -- store, gr0, P2EXPLOSION1POS
  42 => b"00001_0000_10_010000111110", -- store, gr0, P2EXPLOSION1ACTIVE
  43 => b"00001_0000_10_010000111101", -- store, gr0, P2EXPLOSION1TIME
  44 => b"00001_0000_10_010001000101", -- store, gr0, P2EXPLOSION2POS
  45 => b"00001_0000_10_010001000100", -- store, gr0, P2EXPLOSION2ACTIVE
  46 => b"00001_0000_10_010001000011", -- store, gr0, P2EXPLOSION2TIME
  47 => b"00001_0000_10_010001001011", -- store, gr0, P2EXPLOSION3POS
  48 => b"00001_0000_10_010001001010", -- store, gr0, P2EXPLOSION3ACTIVE
  49 => b"00001_0000_10_010001001001", -- store, gr0, P2EXPLOSION3TIME
  50 => b"00000_0000_01_000000000000", -- load, gr0
  51 => b"00000_0000_00_000000000000", -- 0
  52 => b"00000_0011_01_000000000000", -- load, gr3
  53 => b"00000_0000_00_000011000011", -- 195
  54 => b"00001_0000_10_010001010011", -- store, gr0, MOVE
  55 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
  56 => b"00001_0011_10_010001010011", -- store, gr3, MOVE
  57 => b"00011_0010_00_010001010011", -- sub, gr2, MOVE
  58 => b"00110_0000_01_000000000000", -- beq
  59 => b"00000_0000_00_000001000111", -- INITEND
  60 => b"10000_0000_00_000000000000", -- tpoint, gr0
  61 => b"01111_0001_00_000000000000", -- tread, gr1
  62 => b"00011_0001_00_010001010111", -- sub, gr1, WALL
  63 => b"00110_0000_01_000000000000", -- beq
  64 => b"00000_0000_00_000001000011", -- INCREASE
  65 => b"00000_0001_00_010001011000", -- load, gr1, BREAKABLE
  66 => b"01110_0001_00_000000000000", -- twrite, gr1
  67 => b"00010_0000_01_000000000000", -- add, gr0
  68 => b"00000_0000_00_000000000001", -- 1
  69 => b"00100_0000_01_000000000000", -- jump
  70 => b"00000_0000_00_000000110110", -- INITLOOP
  71 => b"00000_0000_00_010001010110", -- load, gr0, GRASS
  72 => b"00000_0001_01_000000000000", -- load, gr1
  73 => b"00000_0000_00_000000010000", -- 16
  74 => b"10000_0001_00_000000000000", -- tpoint, gr1
  75 => b"01110_0000_00_000000000000", -- twrite, gr0
  76 => b"00010_0001_01_000000000000", -- add, gr1
  77 => b"00000_0000_00_000000000001", -- 1
  78 => b"10000_0001_00_000000000000", -- tpoint, gr1
  79 => b"01110_0000_00_000000000000", -- twrite, gr0
  80 => b"00010_0001_01_000000000000", -- add, gr1
  81 => b"00000_0000_00_000000001110", -- 14
  82 => b"10000_0001_00_000000000000", -- tpoint, gr1
  83 => b"01110_0000_00_000000000000", -- twrite, gr0
  84 => b"00000_0001_01_000000000000", -- load, gr1
  85 => b"00000_0000_00_000010110010", -- 178
  86 => b"10000_0001_00_000000000000", -- tpoint, gr1
  87 => b"01110_0000_00_000000000000", -- twrite, gr0
  88 => b"00011_0001_01_000000000000", -- sub, gr1
  89 => b"00000_0000_00_000000000001", -- 1
  90 => b"10000_0001_00_000000000000", -- tpoint, gr1
  91 => b"01110_0000_00_000000000000", -- twrite, gr0
  92 => b"00011_0001_01_000000000000", -- sub, gr1
  93 => b"00000_0000_00_000000001110", -- 14
  94 => b"10000_0001_00_000000000000", -- tpoint, gr1
  95 => b"01110_0000_00_000000000000", -- twrite, gr0
  96 => b"00100_0000_01_000000000000", -- jump
  97 => b"00000_0000_00_000010101000", -- CHECKDEATH
  98 => b"00100_0000_01_000000000000", -- jump
  99 => b"00000_0000_00_000001101110", -- CHECKBOMBDEATH
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_001110000010", -- CONTROL
 102 => b"00100_0000_01_000000000000", -- jump
 103 => b"00000_0000_00_001010111100", -- BUTTON
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000110101101", -- TICKBOMBS
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000011100110", -- TICKEXPLOSIONS
 108 => b"00100_0000_01_000000000000", -- jump
 109 => b"00000_0000_00_000001100000", -- MAIN
 110 => b"00000_0010_01_000000000000", -- load, gr2
 111 => b"00000_0000_00_000000000001", -- 1
 112 => b"00000_0000_00_010000101000", -- load, gr0, P1BOMB1POS
 113 => b"10000_0000_00_000000000000", -- tpoint, gr0
 114 => b"01111_0001_00_000000000000", -- tread, gr1
 115 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 116 => b"00110_0000_01_000000000000", -- beq
 117 => b"00000_0000_00_000010010110", -- P1BOMB1DETONATE
 118 => b"00000_0000_00_010000101110", -- load, gr0, P1BOMB2POS
 119 => b"10000_0000_00_000000000000", -- tpoint, gr0
 120 => b"01111_0001_00_000000000000", -- tread, gr1
 121 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 122 => b"00110_0000_01_000000000000", -- beq
 123 => b"00000_0000_00_000010011001", -- P1BOMB2DETONATE
 124 => b"00000_0000_00_010000110100", -- load, gr0, P1BOMB3POS
 125 => b"10000_0000_00_000000000000", -- tpoint, gr0
 126 => b"01111_0001_00_000000000000", -- tread, gr1
 127 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 128 => b"00110_0000_01_000000000000", -- beq
 129 => b"00000_0000_00_000010011100", -- P1BOMB3DETONATE
 130 => b"00000_0000_00_010000111010", -- load, gr0, P2BOMB1POS
 131 => b"10000_0000_00_000000000000", -- tpoint, gr0
 132 => b"01111_0001_00_000000000000", -- tread, gr1
 133 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 134 => b"00110_0000_01_000000000000", -- beq
 135 => b"00000_0000_00_000010011111", -- P2BOMB1DETONATE
 136 => b"00000_0000_00_010001000000", -- load, gr0, P2BOMB2POS
 137 => b"10000_0000_00_000000000000", -- tpoint, gr0
 138 => b"01111_0001_00_000000000000", -- tread, gr1
 139 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 140 => b"00110_0000_01_000000000000", -- beq
 141 => b"00000_0000_00_000010100010", -- P2BOMB2DETONATE
 142 => b"00000_0000_00_010001000110", -- load, gr0, P2BOMB3POS
 143 => b"10000_0000_00_000000000000", -- tpoint, gr0
 144 => b"01111_0001_00_000000000000", -- tread, gr1
 145 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 146 => b"00110_0000_01_000000000000", -- beq
 147 => b"00000_0000_00_000010100101", -- P2BOMB3DETONATE
 148 => b"00100_0000_01_000000000000", -- jump
 149 => b"00000_0000_00_000001100100", -- CHECKBOMBDEATH_R
 150 => b"00001_0010_10_010000101001", -- store, gr2, P1BOMB1TIME
 151 => b"00100_0000_01_000000000000", -- jump
 152 => b"00000_0000_00_000001110110", -- P1BOMB1DETONATE_R
 153 => b"00001_0010_10_010000101111", -- store, gr2, P1BOMB2TIME
 154 => b"00100_0000_01_000000000000", -- jump
 155 => b"00000_0000_00_000001111100", -- P1BOMB2DETONATE_R
 156 => b"00001_0010_10_010000110101", -- store, gr2, P1BOMB3TIME
 157 => b"00100_0000_01_000000000000", -- jump
 158 => b"00000_0000_00_000010000010", -- P1BOMB3DETONATE_R
 159 => b"00001_0010_10_010000111011", -- store, gr2, P2BOMB1TIME
 160 => b"00100_0000_01_000000000000", -- jump
 161 => b"00000_0000_00_000010001000", -- P2BOMB1DETONATE_R
 162 => b"00001_0010_10_010001000001", -- store, gr2, P2BOMB2TIME
 163 => b"00100_0000_01_000000000000", -- jump
 164 => b"00000_0000_00_000010001110", -- P2BOMB2DETONATE_R
 165 => b"00001_0010_10_010001000111", -- store, gr2, P2BOMB3TIME
 166 => b"00100_0000_01_000000000000", -- jump
 167 => b"00000_0000_00_000010010100", -- P2BOMB3DETONATE_R
 168 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 169 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 170 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 171 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 172 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 173 => b"01000_0000_01_000000000000", -- mul, gr0
 174 => b"00000_0000_00_000000001111", -- 15
 175 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 176 => b"10000_0000_00_000000000000", -- tpoint, gr0
 177 => b"01111_0001_00_000000000000", -- tread, gr1
 178 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 179 => b"00110_0000_01_000000000000", -- beq
 180 => b"00000_0000_00_000011000000", -- P1DEATH
 181 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
 182 => b"01000_0000_01_000000000000", -- mul, gr0
 183 => b"00000_0000_00_000000001111", -- 15
 184 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
 185 => b"10000_0000_00_000000000000", -- tpoint, gr0
 186 => b"01111_0001_00_000000000000", -- tread, gr1
 187 => b"00011_0001_00_010001011001", -- sub, gr1, EXPLOSION
 188 => b"00110_0000_01_000000000000", -- beq
 189 => b"00000_0000_00_000011010011", -- P2DEATH
 190 => b"00100_0000_01_000000000000", -- jump
 191 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 192 => b"00000_0000_01_000000000000", -- load, gr0
 193 => b"00000_0000_00_000000000001", -- 1
 194 => b"00001_0000_10_010000100110", -- store, gr0, P1DEAD
 195 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 196 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 197 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 198 => b"01000_0000_01_000000000000", -- mul, gr0
 199 => b"00000_0000_00_000000001111", -- 15
 200 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 201 => b"10000_0000_00_000000000000", -- tpoint, gr0
 202 => b"00000_0000_01_000000000000", -- load, gr0
 203 => b"00000_0000_00_000000000101", -- 5
 204 => b"01110_0000_00_000000000000", -- twrite, gr0
 205 => b"00000_1100_01_000000000000", -- load, gr12
 206 => b"00000_0000_00_000000000000", -- 0
 207 => b"00000_1101_01_000000000000", -- load, gr13
 208 => b"00000_0000_00_000000010000", -- 16
 209 => b"00100_0000_01_000000000000", -- jump
 210 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 211 => b"00000_0000_01_000000000000", -- load, gr0
 212 => b"00000_0000_00_000000000001", -- 1
 213 => b"00001_0000_10_010000100111", -- store, gr0, P2DEAD
 214 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 215 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 216 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
 217 => b"01000_0000_01_000000000000", -- mul, gr0
 218 => b"00000_0000_00_000000001111", -- 15
 219 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
 220 => b"10000_0000_00_000000000000", -- tpoint, gr0
 221 => b"00000_0000_01_000000000000", -- load, gr0
 222 => b"00000_0000_00_000000000101", -- 5
 223 => b"01110_0000_00_000000000000", -- twrite, gr0
 224 => b"00000_1110_01_000000000000", -- load, gr14
 225 => b"00000_0000_00_000000000000", -- 0
 226 => b"00000_1111_01_000000000000", -- load, gr15
 227 => b"00000_0000_00_000000010000", -- 16
 228 => b"00100_0000_01_000000000000", -- jump
 229 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 230 => b"00000_0000_00_010000101100", -- load, gr0, P1EXPLOSION1ACTIVE
 231 => b"00011_0000_01_000000000000", -- sub, gr0
 232 => b"00000_0000_00_000000000001", -- 1
 233 => b"00111_0000_01_000000000000", -- bne
 234 => b"00000_0000_00_000011110100", -- P1EXPLOSION2
 235 => b"00000_0000_00_010000101011", -- load, gr0, P1EXPLOSION1TIME
 236 => b"00011_0000_01_000000000000", -- sub, gr0
 237 => b"00000_0000_00_000000000001", -- 1
 238 => b"00001_0000_10_010000101011", -- store, gr0, P1EXPLOSION1TIME
 239 => b"00000_0000_01_000000000000", -- load, gr0
 240 => b"00000_0000_00_000000000000", -- 0
 241 => b"00011_0000_00_010000101011", -- sub, gr0, P1EXPLOSION1TIME
 242 => b"00110_0000_01_000000000000", -- beq
 243 => b"00000_0000_00_000100111100", -- P1EXPLOSION1FADE
 244 => b"00000_0000_00_010000110010", -- load, gr0, P1EXPLOSION2ACTIVE
 245 => b"00011_0000_01_000000000000", -- sub, gr0
 246 => b"00000_0000_00_000000000001", -- 1
 247 => b"00111_0000_01_000000000000", -- bne
 248 => b"00000_0000_00_000100000010", -- P1EXPLOSION3
 249 => b"00000_0000_00_010000110001", -- load, gr0, P1EXPLOSION2TIME
 250 => b"00011_0000_01_000000000000", -- sub, gr0
 251 => b"00000_0000_00_000000000001", -- 1
 252 => b"00001_0000_10_010000110001", -- store, gr0, P1EXPLOSION2TIME
 253 => b"00000_0000_01_000000000000", -- load, gr0
 254 => b"00000_0000_00_000000000000", -- 0
 255 => b"00011_0000_00_010000110001", -- sub, gr0, P1EXPLOSION2TIME
 256 => b"00110_0000_01_000000000000", -- beq
 257 => b"00000_0000_00_000101000010", -- P1EXPLOSION2FADE
 258 => b"00000_0000_00_010000111000", -- load, gr0, P1EXPLOSION3ACTIVE
 259 => b"00011_0000_01_000000000000", -- sub, gr0
 260 => b"00000_0000_00_000000000001", -- 1
 261 => b"00111_0000_01_000000000000", -- bne
 262 => b"00000_0000_00_000100010000", -- P2EXPLOSION1
 263 => b"00000_0000_00_010000110111", -- load, gr0, P1EXPLOSION3TIME
 264 => b"00011_0000_01_000000000000", -- sub, gr0
 265 => b"00000_0000_00_000000000001", -- 1
 266 => b"00001_0000_10_010000110111", -- store, gr0, P1EXPLOSION3TIME
 267 => b"00000_0000_01_000000000000", -- load, gr0
 268 => b"00000_0000_00_000000000000", -- 0
 269 => b"00011_0000_00_010000110111", -- sub, gr0, P1EXPLOSION3TIME
 270 => b"00110_0000_01_000000000000", -- beq
 271 => b"00000_0000_00_000101001000", -- P1EXPLOSION3FADE
 272 => b"00000_0000_00_010000111110", -- load, gr0, P2EXPLOSION1ACTIVE
 273 => b"00011_0000_01_000000000000", -- sub, gr0
 274 => b"00000_0000_00_000000000001", -- 1
 275 => b"00111_0000_01_000000000000", -- bne
 276 => b"00000_0000_00_000100011110", -- P2EXPLOSION2
 277 => b"00000_0000_00_010000111101", -- load, gr0, P2EXPLOSION1TIME
 278 => b"00011_0000_01_000000000000", -- sub, gr0
 279 => b"00000_0000_00_000000000001", -- 1
 280 => b"00001_0000_10_010000111101", -- store, gr0, P2EXPLOSION1TIME
 281 => b"00000_0000_01_000000000000", -- load, gr0
 282 => b"00000_0000_00_000000000000", -- 0
 283 => b"00011_0000_00_010000111101", -- sub, gr0, P2EXPLOSION1TIME
 284 => b"00110_0000_01_000000000000", -- beq
 285 => b"00000_0000_00_000101001110", -- P2EXPLOSION1FADE
 286 => b"00000_0000_00_010001000100", -- load, gr0, P2EXPLOSION2ACTIVE
 287 => b"00011_0000_01_000000000000", -- sub, gr0
 288 => b"00000_0000_00_000000000001", -- 1
 289 => b"00111_0000_01_000000000000", -- bne
 290 => b"00000_0000_00_000100101100", -- P2EXPLOSION3
 291 => b"00000_0000_00_010001000011", -- load, gr0, P2EXPLOSION2TIME
 292 => b"00011_0000_01_000000000000", -- sub, gr0
 293 => b"00000_0000_00_000000000001", -- 1
 294 => b"00001_0000_10_010001000011", -- store, gr0, P2EXPLOSION2TIME
 295 => b"00000_0000_01_000000000000", -- load, gr0
 296 => b"00000_0000_00_000000000000", -- 0
 297 => b"00011_0000_00_010001000011", -- sub, gr0, P2EXPLOSION2TIME
 298 => b"00110_0000_01_000000000000", -- beq
 299 => b"00000_0000_00_000101010100", -- P2EXPLOSION2FADE
 300 => b"00000_0000_00_010001001010", -- load, gr0, P2EXPLOSION3ACTIVE
 301 => b"00011_0000_01_000000000000", -- sub, gr0
 302 => b"00000_0000_00_000000000001", -- 1
 303 => b"00111_0000_01_000000000000", -- bne
 304 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 305 => b"00000_0000_00_010001001001", -- load, gr0, P2EXPLOSION3TIME
 306 => b"00011_0000_01_000000000000", -- sub, gr0
 307 => b"00000_0000_00_000000000001", -- 1
 308 => b"00001_0000_10_010001001001", -- store, gr0, P2EXPLOSION3TIME
 309 => b"00000_0000_01_000000000000", -- load, gr0
 310 => b"00000_0000_00_000000000000", -- 0
 311 => b"00011_0000_00_010001001001", -- sub, gr0, P2EXPLOSION3TIME
 312 => b"00110_0000_01_000000000000", -- beq
 313 => b"00000_0000_00_000101011010", -- P2EXPLOSION3FADE
 314 => b"00100_0000_01_000000000000", -- jump
 315 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 316 => b"00000_0000_01_000000000000", -- load, gr0
 317 => b"00000_0000_00_000000000000", -- 0
 318 => b"00001_0000_10_010000101100", -- store, gr0, P1EXPLOSION1ACTIVE
 319 => b"00000_0100_00_010000101101", -- load, gr4, P1EXPLOSION1POS
 320 => b"00100_0000_01_000000000000", -- jump
 321 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 322 => b"00000_0000_01_000000000000", -- load, gr0
 323 => b"00000_0000_00_000000000000", -- 0
 324 => b"00001_0000_10_010000110010", -- store, gr0, P1EXPLOSION2ACTIVE
 325 => b"00000_0100_00_010000110011", -- load, gr4, P1EXPLOSION2POS
 326 => b"00100_0000_01_000000000000", -- jump
 327 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 328 => b"00000_0000_01_000000000000", -- load, gr0
 329 => b"00000_0000_00_000000000000", -- 0
 330 => b"00001_0000_10_010000111000", -- store, gr0, P1EXPLOSION3ACTIVE
 331 => b"00000_0100_00_010000111001", -- load, gr4, P1EXPLOSION3POS
 332 => b"00100_0000_01_000000000000", -- jump
 333 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 334 => b"00000_0000_01_000000000000", -- load, gr0
 335 => b"00000_0000_00_000000000000", -- 0
 336 => b"00001_0000_10_010000111110", -- store, gr0, P2EXPLOSION1ACTIVE
 337 => b"00000_0100_00_010000111111", -- load, gr4, P2EXPLOSION1POS
 338 => b"00100_0000_01_000000000000", -- jump
 339 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 340 => b"00000_0000_01_000000000000", -- load, gr0
 341 => b"00000_0000_00_000000000000", -- 0
 342 => b"00001_0000_10_010001000100", -- store, gr0, P2EXPLOSION2ACTIVE
 343 => b"00000_0100_00_010001000101", -- load, gr4, P2EXPLOSION2POS
 344 => b"00100_0000_01_000000000000", -- jump
 345 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 346 => b"00000_0000_01_000000000000", -- load, gr0
 347 => b"00000_0000_00_000000000000", -- 0
 348 => b"00001_0000_10_010001001010", -- store, gr0, P2EXPLOSION3ACTIVE
 349 => b"00000_0100_00_010001001011", -- load, gr4, P2EXPLOSION3POS
 350 => b"00100_0000_01_000000000000", -- jump
 351 => b"00000_0000_00_000101100000", -- FADEEXPLOSION
 352 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 353 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 354 => b"00000_0011_00_010001010110", -- load, gr3, GRASS
 355 => b"10000_0010_00_000000000000", -- tpoint, gr2
 356 => b"01110_0011_00_000000000000", -- twrite, gr3
 357 => b"00010_0010_01_000000000000", -- add, gr2
 358 => b"00000_0000_00_000000000001", -- 1
 359 => b"10000_0010_00_000000000000", -- tpoint, gr2
 360 => b"01111_0000_00_000000000000", -- tread, gr0
 361 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 362 => b"00110_0000_01_000000000000", -- beq
 363 => b"00000_0000_00_000101110101", -- FADELEFT
 364 => b"01110_0011_00_000000000000", -- twrite, gr3
 365 => b"00010_0010_01_000000000000", -- add, gr2
 366 => b"00000_0000_00_000000000001", -- 1
 367 => b"10000_0010_00_000000000000", -- tpoint, gr2
 368 => b"01111_0000_00_000000000000", -- tread, gr0
 369 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 370 => b"00110_0000_01_000000000000", -- beq
 371 => b"00000_0000_00_000101110101", -- FADELEFT
 372 => b"01110_0011_00_000000000000", -- twrite, gr3
 373 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 374 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 375 => b"00011_0010_01_000000000000", -- sub, gr2
 376 => b"00000_0000_00_000000000001", -- 1
 377 => b"10000_0010_00_000000000000", -- tpoint, gr2
 378 => b"01111_0000_00_000000000000", -- tread, gr0
 379 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 380 => b"00110_0000_01_000000000000", -- beq
 381 => b"00000_0000_00_000110000111", -- FADEDOWN
 382 => b"01110_0011_00_000000000000", -- twrite, gr3
 383 => b"00011_0010_01_000000000000", -- sub, gr2
 384 => b"00000_0000_00_000000000001", -- 1
 385 => b"10000_0010_00_000000000000", -- tpoint, gr2
 386 => b"01111_0000_00_000000000000", -- tread, gr0
 387 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 388 => b"00110_0000_01_000000000000", -- beq
 389 => b"00000_0000_00_000110000111", -- FADEDOWN
 390 => b"01110_0011_00_000000000000", -- twrite, gr3
 391 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 392 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 393 => b"00010_0010_01_000000000000", -- add, gr2
 394 => b"00000_0000_00_000000001111", -- 15
 395 => b"10000_0010_00_000000000000", -- tpoint, gr2
 396 => b"01111_0000_00_000000000000", -- tread, gr0
 397 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 398 => b"00110_0000_01_000000000000", -- beq
 399 => b"00000_0000_00_000110011001", -- FADEUP
 400 => b"01110_0011_00_000000000000", -- twrite, gr3
 401 => b"00010_0010_01_000000000000", -- add, gr2
 402 => b"00000_0000_00_000000001111", -- 15
 403 => b"10000_0010_00_000000000000", -- tpoint, gr2
 404 => b"01111_0000_00_000000000000", -- tread, gr0
 405 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 406 => b"00110_0000_01_000000000000", -- beq
 407 => b"00000_0000_00_000110011001", -- FADEUP
 408 => b"01110_0011_00_000000000000", -- twrite, gr3
 409 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 410 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 411 => b"00011_0010_01_000000000000", -- sub, gr2
 412 => b"00000_0000_00_000000001111", -- 15
 413 => b"10000_0010_00_000000000000", -- tpoint, gr2
 414 => b"01111_0000_00_000000000000", -- tread, gr0
 415 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 416 => b"00110_0000_01_000000000000", -- beq
 417 => b"00000_0000_00_000011100110", -- TICKEXPLOSIONS
 418 => b"01110_0011_00_000000000000", -- twrite, gr3
 419 => b"00011_0010_01_000000000000", -- sub, gr2
 420 => b"00000_0000_00_000000001111", -- 15
 421 => b"10000_0010_00_000000000000", -- tpoint, gr2
 422 => b"01111_0000_00_000000000000", -- tread, gr0
 423 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 424 => b"00110_0000_01_000000000000", -- beq
 425 => b"00000_0000_00_000011100110", -- TICKEXPLOSIONS
 426 => b"01110_0011_00_000000000000", -- twrite, gr3
 427 => b"00100_0000_01_000000000000", -- jump
 428 => b"00000_0000_00_000011100110", -- TICKEXPLOSIONS
 429 => b"00000_0000_00_010000101010", -- load, gr0, P1BOMB1ACTIVE
 430 => b"00011_0000_01_000000000000", -- sub, gr0
 431 => b"00000_0000_00_000000000001", -- 1
 432 => b"00111_0000_01_000000000000", -- bne
 433 => b"00000_0000_00_000110111011", -- P1BOMB2
 434 => b"00000_0000_00_010000101001", -- load, gr0, P1BOMB1TIME
 435 => b"00011_0000_01_000000000000", -- sub, gr0
 436 => b"00000_0000_00_000000000001", -- 1
 437 => b"00001_0000_10_010000101001", -- store, gr0, P1BOMB1TIME
 438 => b"00000_0000_01_000000000000", -- load, gr0
 439 => b"00000_0000_00_000000000000", -- 0
 440 => b"00011_0000_00_010000101001", -- sub, gr0, P1BOMB1TIME
 441 => b"00110_0000_01_000000000000", -- beq
 442 => b"00000_0000_00_001000000011", -- P1EXPLOSION1INIT
 443 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMB2ACTIVE
 444 => b"00011_0000_01_000000000000", -- sub, gr0
 445 => b"00000_0000_00_000000000001", -- 1
 446 => b"00111_0000_01_000000000000", -- bne
 447 => b"00000_0000_00_000111001001", -- P1BOMB3
 448 => b"00000_0000_00_010000101111", -- load, gr0, P1BOMB2TIME
 449 => b"00011_0000_01_000000000000", -- sub, gr0
 450 => b"00000_0000_00_000000000001", -- 1
 451 => b"00001_0000_10_010000101111", -- store, gr0, P1BOMB2TIME
 452 => b"00000_0000_01_000000000000", -- load, gr0
 453 => b"00000_0000_00_000000000000", -- 0
 454 => b"00011_0000_00_010000101111", -- sub, gr0, P1BOMB2TIME
 455 => b"00110_0000_01_000000000000", -- beq
 456 => b"00000_0000_00_001000010101", -- P1EXPLOSION2INIT
 457 => b"00000_0000_00_010000110110", -- load, gr0, P1BOMB3ACTIVE
 458 => b"00011_0000_01_000000000000", -- sub, gr0
 459 => b"00000_0000_00_000000000001", -- 1
 460 => b"00111_0000_01_000000000000", -- bne
 461 => b"00000_0000_00_000111010111", -- P2BOMB1
 462 => b"00000_0000_00_010000110101", -- load, gr0, P1BOMB3TIME
 463 => b"00011_0000_01_000000000000", -- sub, gr0
 464 => b"00000_0000_00_000000000001", -- 1
 465 => b"00001_0000_10_010000110101", -- store, gr0, P1BOMB3TIME
 466 => b"00000_0000_01_000000000000", -- load, gr0
 467 => b"00000_0000_00_000000000000", -- 0
 468 => b"00011_0000_00_010000110101", -- sub, gr0, P1BOMB3TIME
 469 => b"00110_0000_01_000000000000", -- beq
 470 => b"00000_0000_00_001000100111", -- P1EXPLOSION3INIT
 471 => b"00000_0000_00_010000111100", -- load, gr0, P2BOMB1ACTIVE
 472 => b"00011_0000_01_000000000000", -- sub, gr0
 473 => b"00000_0000_00_000000000001", -- 1
 474 => b"00111_0000_01_000000000000", -- bne
 475 => b"00000_0000_00_000111100101", -- P2BOMB2
 476 => b"00000_0000_00_010000111011", -- load, gr0, P2BOMB1TIME
 477 => b"00011_0000_01_000000000000", -- sub, gr0
 478 => b"00000_0000_00_000000000001", -- 1
 479 => b"00001_0000_10_010000111011", -- store, gr0, P2BOMB1TIME
 480 => b"00000_0000_01_000000000000", -- load, gr0
 481 => b"00000_0000_00_000000000000", -- 0
 482 => b"00011_0000_00_010000111011", -- sub, gr0, P2BOMB1TIME
 483 => b"00110_0000_01_000000000000", -- beq
 484 => b"00000_0000_00_001000111001", -- P2EXPLOSION1INIT
 485 => b"00000_0000_00_010001000010", -- load, gr0, P2BOMB2ACTIVE
 486 => b"00011_0000_01_000000000000", -- sub, gr0
 487 => b"00000_0000_00_000000000001", -- 1
 488 => b"00111_0000_01_000000000000", -- bne
 489 => b"00000_0000_00_000111110011", -- P2BOMB3
 490 => b"00000_0000_00_010001000001", -- load, gr0, P2BOMB2TIME
 491 => b"00011_0000_01_000000000000", -- sub, gr0
 492 => b"00000_0000_00_000000000001", -- 1
 493 => b"00001_0000_10_010001000001", -- store, gr0, P2BOMB2TIME
 494 => b"00000_0000_01_000000000000", -- load, gr0
 495 => b"00000_0000_00_000000000000", -- 0
 496 => b"00011_0000_00_010001000001", -- sub, gr0, P2BOMB2TIME
 497 => b"00110_0000_01_000000000000", -- beq
 498 => b"00000_0000_00_001001001011", -- P2EXPLOSION2INIT
 499 => b"00000_0000_00_010001001000", -- load, gr0, P2BOMB3ACTIVE
 500 => b"00011_0000_01_000000000000", -- sub, gr0
 501 => b"00000_0000_00_000000000001", -- 1
 502 => b"00111_0000_01_000000000000", -- bne
 503 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 504 => b"00000_0000_00_010001000111", -- load, gr0, P2BOMB3TIME
 505 => b"00011_0000_01_000000000000", -- sub, gr0
 506 => b"00000_0000_00_000000000001", -- 1
 507 => b"00001_0000_10_010001000111", -- store, gr0, P2BOMB3TIME
 508 => b"00000_0000_01_000000000000", -- load, gr0
 509 => b"00000_0000_00_000000000000", -- 0
 510 => b"00011_0000_00_010001000111", -- sub, gr0, P2BOMB3TIME
 511 => b"00110_0000_01_000000000000", -- beq
 512 => b"00000_0000_00_001001011101", -- P2EXPLOSION3INIT
 513 => b"00100_0000_01_000000000000", -- jump
 514 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 515 => b"00000_0000_01_000000000000", -- load, gr0
 516 => b"00000_0000_00_000000000000", -- 0
 517 => b"00001_0000_10_010000101010", -- store, gr0, P1BOMB1ACTIVE
 518 => b"00000_0000_00_010000101000", -- load, gr0, P1BOMB1POS
 519 => b"00001_0000_10_010000101101", -- store, gr0, P1EXPLOSION1POS
 520 => b"00000_0000_01_000000000000", -- load, gr0
 521 => b"00000_0000_00_000000000001", -- 1
 522 => b"00001_0000_10_010000101100", -- store, gr0, P1EXPLOSION1ACTIVE
 523 => b"00000_0000_01_000000000000", -- load, gr0
 524 => b"00000_0000_00_000000000010", -- 2
 525 => b"00001_0000_10_010000101011", -- store, gr0, P1EXPLOSION1TIME
 526 => b"00000_0000_00_010001001100", -- load, gr0, P1BOMBCOUNT
 527 => b"00011_0000_01_000000000000", -- sub, gr0
 528 => b"00000_0000_00_000000000001", -- 1
 529 => b"00001_0000_10_010001001100", -- store, gr0, P1BOMBCOUNT
 530 => b"00000_0100_00_010000101000", -- load, gr4, P1BOMB1POS
 531 => b"00100_0000_01_000000000000", -- jump
 532 => b"00000_0000_00_001001101111", -- EXPLODE
 533 => b"00000_0000_01_000000000000", -- load, gr0
 534 => b"00000_0000_00_000000000000", -- 0
 535 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMB2ACTIVE
 536 => b"00000_0000_00_010000101110", -- load, gr0, P1BOMB2POS
 537 => b"00001_0000_10_010000110011", -- store, gr0, P1EXPLOSION2POS
 538 => b"00000_0000_01_000000000000", -- load, gr0
 539 => b"00000_0000_00_000000000001", -- 1
 540 => b"00001_0000_10_010000110010", -- store, gr0, P1EXPLOSION2ACTIVE
 541 => b"00000_0000_01_000000000000", -- load, gr0
 542 => b"00000_0000_00_000000000010", -- 2
 543 => b"00001_0000_10_010000110001", -- store, gr0, P1EXPLOSION2TIME
 544 => b"00000_0000_00_010001001100", -- load, gr0, P1BOMBCOUNT
 545 => b"00011_0000_01_000000000000", -- sub, gr0
 546 => b"00000_0000_00_000000000001", -- 1
 547 => b"00001_0000_10_010001001100", -- store, gr0, P1BOMBCOUNT
 548 => b"00000_0100_00_010000101110", -- load, gr4, P1BOMB2POS
 549 => b"00100_0000_01_000000000000", -- jump
 550 => b"00000_0000_00_001001101111", -- EXPLODE
 551 => b"00000_0000_01_000000000000", -- load, gr0
 552 => b"00000_0000_00_000000000000", -- 0
 553 => b"00001_0000_10_010000110110", -- store, gr0, P1BOMB3ACTIVE
 554 => b"00000_0000_00_010000110100", -- load, gr0, P1BOMB3POS
 555 => b"00001_0000_10_010000111001", -- store, gr0, P1EXPLOSION3POS
 556 => b"00000_0000_01_000000000000", -- load, gr0
 557 => b"00000_0000_00_000000000001", -- 1
 558 => b"00001_0000_10_010000111000", -- store, gr0, P1EXPLOSION3ACTIVE
 559 => b"00000_0000_01_000000000000", -- load, gr0
 560 => b"00000_0000_00_000000000010", -- 2
 561 => b"00001_0000_10_010000110111", -- store, gr0, P1EXPLOSION3TIME
 562 => b"00000_0000_00_010001001100", -- load, gr0, P1BOMBCOUNT
 563 => b"00011_0000_01_000000000000", -- sub, gr0
 564 => b"00000_0000_00_000000000001", -- 1
 565 => b"00001_0000_10_010001001100", -- store, gr0, P1BOMBCOUNT
 566 => b"00000_0100_00_010000110100", -- load, gr4, P1BOMB3POS
 567 => b"00100_0000_01_000000000000", -- jump
 568 => b"00000_0000_00_001001101111", -- EXPLODE
 569 => b"00000_0000_01_000000000000", -- load, gr0
 570 => b"00000_0000_00_000000000000", -- 0
 571 => b"00001_0000_10_010000111100", -- store, gr0, P2BOMB1ACTIVE
 572 => b"00000_0000_00_010000111010", -- load, gr0, P2BOMB1POS
 573 => b"00001_0000_10_010000111111", -- store, gr0, P2EXPLOSION1POS
 574 => b"00000_0000_01_000000000000", -- load, gr0
 575 => b"00000_0000_00_000000000001", -- 1
 576 => b"00001_0000_10_010000111110", -- store, gr0, P2EXPLOSION1ACTIVE
 577 => b"00000_0000_01_000000000000", -- load, gr0
 578 => b"00000_0000_00_000000000010", -- 2
 579 => b"00001_0000_10_010000111101", -- store, gr0, P2EXPLOSION1TIME
 580 => b"00000_0000_00_010001001101", -- load, gr0, P2BOMBCOUNT
 581 => b"00011_0000_01_000000000000", -- sub, gr0
 582 => b"00000_0000_00_000000000001", -- 1
 583 => b"00001_0000_10_010001001101", -- store, gr0, P2BOMBCOUNT
 584 => b"00000_0100_00_010000111010", -- load, gr4, P2BOMB1POS
 585 => b"00100_0000_01_000000000000", -- jump
 586 => b"00000_0000_00_001001101111", -- EXPLODE
 587 => b"00000_0000_01_000000000000", -- load, gr0
 588 => b"00000_0000_00_000000000000", -- 0
 589 => b"00001_0000_10_010001000010", -- store, gr0, P2BOMB2ACTIVE
 590 => b"00000_0000_00_010001000000", -- load, gr0, P2BOMB2POS
 591 => b"00001_0000_10_010001000101", -- store, gr0, P2EXPLOSION2POS
 592 => b"00000_0000_01_000000000000", -- load, gr0
 593 => b"00000_0000_00_000000000001", -- 1
 594 => b"00001_0000_10_010001000100", -- store, gr0, P2EXPLOSION2ACTIVE
 595 => b"00000_0000_01_000000000000", -- load, gr0
 596 => b"00000_0000_00_000000000010", -- 2
 597 => b"00001_0000_10_010001000011", -- store, gr0, P2EXPLOSION2TIME
 598 => b"00000_0000_00_010001001101", -- load, gr0, P2BOMBCOUNT
 599 => b"00011_0000_01_000000000000", -- sub, gr0
 600 => b"00000_0000_00_000000000001", -- 1
 601 => b"00001_0000_10_010001001101", -- store, gr0, P2BOMBCOUNT
 602 => b"00000_0100_00_010001000000", -- load, gr4, P2BOMB2POS
 603 => b"00100_0000_01_000000000000", -- jump
 604 => b"00000_0000_00_001001101111", -- EXPLODE
 605 => b"00000_0000_01_000000000000", -- load, gr0
 606 => b"00000_0000_00_000000000000", -- 0
 607 => b"00001_0000_10_010001001000", -- store, gr0, P2BOMB3ACTIVE
 608 => b"00000_0000_00_010001000110", -- load, gr0, P2BOMB3POS
 609 => b"00001_0000_10_010001001011", -- store, gr0, P2EXPLOSION3POS
 610 => b"00000_0000_01_000000000000", -- load, gr0
 611 => b"00000_0000_00_000000000001", -- 1
 612 => b"00001_0000_10_010001001010", -- store, gr0, P2EXPLOSION3ACTIVE
 613 => b"00000_0000_01_000000000000", -- load, gr0
 614 => b"00000_0000_00_000000000010", -- 2
 615 => b"00001_0000_10_010001001001", -- store, gr0, P2EXPLOSION3TIME
 616 => b"00000_0000_00_010001001101", -- load, gr0, P2BOMBCOUNT
 617 => b"00011_0000_01_000000000000", -- sub, gr0
 618 => b"00000_0000_00_000000000001", -- 1
 619 => b"00001_0000_10_010001001101", -- store, gr0, P2BOMBCOUNT
 620 => b"00000_0100_00_010001000110", -- load, gr4, P2BOMB3POS
 621 => b"00100_0000_01_000000000000", -- jump
 622 => b"00000_0000_00_001001101111", -- EXPLODE
 623 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 624 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 625 => b"00000_0011_00_010001011001", -- load, gr3, EXPLOSION
 626 => b"10000_0010_00_000000000000", -- tpoint, gr2
 627 => b"01110_0011_00_000000000000", -- twrite, gr3
 628 => b"00010_0010_01_000000000000", -- add, gr2
 629 => b"00000_0000_00_000000000001", -- 1
 630 => b"10000_0010_00_000000000000", -- tpoint, gr2
 631 => b"01111_0000_00_000000000000", -- tread, gr0
 632 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 633 => b"00110_0000_01_000000000000", -- beq
 634 => b"00000_0000_00_001010000100", -- EXPLODELEFT
 635 => b"01110_0011_00_000000000000", -- twrite, gr3
 636 => b"00010_0010_01_000000000000", -- add, gr2
 637 => b"00000_0000_00_000000000001", -- 1
 638 => b"10000_0010_00_000000000000", -- tpoint, gr2
 639 => b"01111_0000_00_000000000000", -- tread, gr0
 640 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 641 => b"00110_0000_01_000000000000", -- beq
 642 => b"00000_0000_00_001010000100", -- EXPLODELEFT
 643 => b"01110_0011_00_000000000000", -- twrite, gr3
 644 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 645 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 646 => b"00011_0010_01_000000000000", -- sub, gr2
 647 => b"00000_0000_00_000000000001", -- 1
 648 => b"10000_0010_00_000000000000", -- tpoint, gr2
 649 => b"01111_0000_00_000000000000", -- tread, gr0
 650 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 651 => b"00110_0000_01_000000000000", -- beq
 652 => b"00000_0000_00_001010010110", -- EXPLODEDOWN
 653 => b"01110_0011_00_000000000000", -- twrite, gr3
 654 => b"00011_0010_01_000000000000", -- sub, gr2
 655 => b"00000_0000_00_000000000001", -- 1
 656 => b"10000_0010_00_000000000000", -- tpoint, gr2
 657 => b"01111_0000_00_000000000000", -- tread, gr0
 658 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 659 => b"00110_0000_01_000000000000", -- beq
 660 => b"00000_0000_00_001010010110", -- EXPLODEDOWN
 661 => b"01110_0011_00_000000000000", -- twrite, gr3
 662 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 663 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 664 => b"00010_0010_01_000000000000", -- add, gr2
 665 => b"00000_0000_00_000000001111", -- 15
 666 => b"10000_0010_00_000000000000", -- tpoint, gr2
 667 => b"01111_0000_00_000000000000", -- tread, gr0
 668 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 669 => b"00110_0000_01_000000000000", -- beq
 670 => b"00000_0000_00_001010101000", -- EXPLODEUP
 671 => b"01110_0011_00_000000000000", -- twrite, gr3
 672 => b"00010_0010_01_000000000000", -- add, gr2
 673 => b"00000_0000_00_000000001111", -- 15
 674 => b"10000_0010_00_000000000000", -- tpoint, gr2
 675 => b"01111_0000_00_000000000000", -- tread, gr0
 676 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 677 => b"00110_0000_01_000000000000", -- beq
 678 => b"00000_0000_00_001010101000", -- EXPLODEUP
 679 => b"01110_0011_00_000000000000", -- twrite, gr3
 680 => b"00001_0100_10_010001010011", -- store, gr4, MOVE
 681 => b"00000_0010_00_010001010011", -- load, gr2, MOVE
 682 => b"00011_0010_01_000000000000", -- sub, gr2
 683 => b"00000_0000_00_000000001111", -- 15
 684 => b"10000_0010_00_000000000000", -- tpoint, gr2
 685 => b"01111_0000_00_000000000000", -- tread, gr0
 686 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 687 => b"00110_0000_01_000000000000", -- beq
 688 => b"00000_0000_00_000110101101", -- TICKBOMBS
 689 => b"01110_0011_00_000000000000", -- twrite, gr3
 690 => b"00011_0010_01_000000000000", -- sub, gr2
 691 => b"00000_0000_00_000000001111", -- 15
 692 => b"10000_0010_00_000000000000", -- tpoint, gr2
 693 => b"01111_0000_00_000000000000", -- tread, gr0
 694 => b"00011_0000_00_010001010111", -- sub, gr0, WALL
 695 => b"00110_0000_01_000000000000", -- beq
 696 => b"00000_0000_00_000110101101", -- TICKBOMBS
 697 => b"01110_0011_00_000000000000", -- twrite, gr3
 698 => b"00100_0000_01_000000000000", -- jump
 699 => b"00000_0000_00_000110101101", -- TICKBOMBS
 700 => b"10101_0000_01_000000000000", -- btn1
 701 => b"00000_0000_00_001011000010", -- BTN1
 702 => b"11010_0000_01_000000000000", -- btn2
 703 => b"00000_0000_00_001100100011", -- BTN2
 704 => b"00100_0000_01_000000000000", -- jump
 705 => b"00000_0000_00_000001101000", -- BUTTON_R
 706 => b"00000_0000_00_010000100110", -- load, gr0, P1DEAD
 707 => b"00011_0000_01_000000000000", -- sub, gr0
 708 => b"00000_0000_00_000000000001", -- 1
 709 => b"00110_0000_01_000000000000", -- beq
 710 => b"00000_0000_00_000000000000", -- INIT
 711 => b"00000_0000_00_010001001100", -- load, gr0, P1BOMBCOUNT
 712 => b"00011_0000_00_010001001110", -- sub, gr0, MAXBOMBS
 713 => b"00110_0000_01_000000000000", -- beq
 714 => b"00000_0000_00_001010111110", -- BTN1_R
 715 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 716 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 717 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 718 => b"01000_0000_01_000000000000", -- mul, gr0
 719 => b"00000_0000_00_000000001111", -- 15
 720 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 721 => b"10000_0000_00_000000000000", -- tpoint, gr0
 722 => b"01111_0001_00_000000000000", -- tread, gr1
 723 => b"00011_0001_00_010001011010", -- sub, gr1, EGG
 724 => b"00110_0000_01_000000000000", -- beq
 725 => b"00000_0000_00_001010111110", -- BTN1_R
 726 => b"00000_0000_00_010000101010", -- load, gr0, P1BOMB1ACTIVE
 727 => b"00011_0000_01_000000000000", -- sub, gr0
 728 => b"00000_0000_00_000000000000", -- 0
 729 => b"00110_0000_01_000000000000", -- beq
 730 => b"00000_0000_00_001011101101", -- P1PLACEBOMB1
 731 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMB2ACTIVE
 732 => b"00011_0000_01_000000000000", -- sub, gr0
 733 => b"00000_0000_00_000000000000", -- 0
 734 => b"00110_0000_01_000000000000", -- beq
 735 => b"00000_0000_00_001011111111", -- P1PLACEBOMB2
 736 => b"00000_0000_00_010000110110", -- load, gr0, P1BOMB3ACTIVE
 737 => b"00011_0000_01_000000000000", -- sub, gr0
 738 => b"00000_0000_00_000000000000", -- 0
 739 => b"00110_0000_01_000000000000", -- beq
 740 => b"00000_0000_00_001100010001", -- P1PLACEBOMB3
 741 => b"00100_0000_01_000000000000", -- jump
 742 => b"00000_0000_00_001010111110", -- BTN1_R
 743 => b"00000_0000_00_010001001100", -- load, gr0, P1BOMBCOUNT
 744 => b"00010_0000_01_000000000000", -- add, gr0
 745 => b"00000_0000_00_000000000001", -- 1
 746 => b"00001_0000_10_010001001100", -- store, gr0, P1BOMBCOUNT
 747 => b"00100_0000_01_000000000000", -- jump
 748 => b"00000_0000_00_001010111110", -- BTN1_R
 749 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 750 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 751 => b"00000_0011_00_010001010000", -- load, gr3, YPOS1
 752 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 753 => b"01000_0011_01_000000000000", -- mul, gr3
 754 => b"00000_0000_00_000000001111", -- 15
 755 => b"00010_0011_00_010001001111", -- add, gr3, XPOS1
 756 => b"10000_0011_00_000000000000", -- tpoint, gr3
 757 => b"01110_0010_00_000000000000", -- twrite, gr2
 758 => b"00000_0000_01_000000000000", -- load, gr0
 759 => b"00000_0000_00_000000000001", -- 1
 760 => b"00001_0000_10_010000101010", -- store, gr0, P1BOMB1ACTIVE
 761 => b"00001_0011_10_010000101000", -- store, gr3, P1BOMB1POS
 762 => b"00000_0000_01_000000000000", -- load, gr0
 763 => b"00000_0000_00_000000010000", -- 16
 764 => b"00001_0000_10_010000101001", -- store, gr0, P1BOMB1TIME
 765 => b"00100_0000_01_000000000000", -- jump
 766 => b"00000_0000_00_001011100111", -- P1INCREASEBOMBCOUNTER
 767 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 768 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 769 => b"00000_0011_00_010001010000", -- load, gr3, YPOS1
 770 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 771 => b"01000_0011_01_000000000000", -- mul, gr3
 772 => b"00000_0000_00_000000001111", -- 15
 773 => b"00010_0011_00_010001001111", -- add, gr3, XPOS1
 774 => b"10000_0011_00_000000000000", -- tpoint, gr3
 775 => b"01110_0010_00_000000000000", -- twrite, gr2
 776 => b"00000_0000_01_000000000000", -- load, gr0
 777 => b"00000_0000_00_000000000001", -- 1
 778 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMB2ACTIVE
 779 => b"00001_0011_10_010000101110", -- store, gr3, P1BOMB2POS
 780 => b"00000_0000_01_000000000000", -- load, gr0
 781 => b"00000_0000_00_000000010000", -- 16
 782 => b"00001_0000_10_010000101111", -- store, gr0, P1BOMB2TIME
 783 => b"00100_0000_01_000000000000", -- jump
 784 => b"00000_0000_00_001011100111", -- P1INCREASEBOMBCOUNTER
 785 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 786 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 787 => b"00000_0011_00_010001010000", -- load, gr3, YPOS1
 788 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 789 => b"01000_0011_01_000000000000", -- mul, gr3
 790 => b"00000_0000_00_000000001111", -- 15
 791 => b"00010_0011_00_010001001111", -- add, gr3, XPOS1
 792 => b"10000_0011_00_000000000000", -- tpoint, gr3
 793 => b"01110_0010_00_000000000000", -- twrite, gr2
 794 => b"00000_0000_01_000000000000", -- load, gr0
 795 => b"00000_0000_00_000000000001", -- 1
 796 => b"00001_0000_10_010000110110", -- store, gr0, P1BOMB3ACTIVE
 797 => b"00001_0011_10_010000110100", -- store, gr3, P1BOMB3POS
 798 => b"00000_0000_01_000000000000", -- load, gr0
 799 => b"00000_0000_00_000000010000", -- 16
 800 => b"00001_0000_10_010000110101", -- store, gr0, P1BOMB3TIME
 801 => b"00100_0000_01_000000000000", -- jump
 802 => b"00000_0000_00_001011100111", -- P1INCREASEBOMBCOUNTER
 803 => b"00000_0000_00_010000100111", -- load, gr0, P2DEAD
 804 => b"00011_0000_01_000000000000", -- sub, gr0
 805 => b"00000_0000_00_000000000001", -- 1
 806 => b"00110_0000_01_000000000000", -- beq
 807 => b"00000_0000_00_000000000000", -- INIT
 808 => b"00000_0000_00_010001001101", -- load, gr0, P2BOMBCOUNT
 809 => b"00011_0000_00_010001001110", -- sub, gr0, MAXBOMBS
 810 => b"00110_0000_01_000000000000", -- beq
 811 => b"00000_0000_00_001011000000", -- BTN2_R
 812 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 813 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 814 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
 815 => b"01000_0000_01_000000000000", -- mul, gr0
 816 => b"00000_0000_00_000000001111", -- 15
 817 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
 818 => b"10000_0000_00_000000000000", -- tpoint, gr0
 819 => b"01111_0001_00_000000000000", -- tread, gr1
 820 => b"00011_0001_00_010001011010", -- sub, gr1, EGG
 821 => b"00110_0000_01_000000000000", -- beq
 822 => b"00000_0000_00_001011000000", -- BTN2_R
 823 => b"00000_0000_00_010000111100", -- load, gr0, P2BOMB1ACTIVE
 824 => b"00011_0000_01_000000000000", -- sub, gr0
 825 => b"00000_0000_00_000000000000", -- 0
 826 => b"00110_0000_01_000000000000", -- beq
 827 => b"00000_0000_00_001101001100", -- P2PLACEBOMB1
 828 => b"00000_0000_00_010001000010", -- load, gr0, P2BOMB2ACTIVE
 829 => b"00011_0000_01_000000000000", -- sub, gr0
 830 => b"00000_0000_00_000000000000", -- 0
 831 => b"00110_0000_01_000000000000", -- beq
 832 => b"00000_0000_00_001101011110", -- P2PLACEBOMB2
 833 => b"00000_0000_00_010001001000", -- load, gr0, P2BOMB3ACTIVE
 834 => b"00011_0000_01_000000000000", -- sub, gr0
 835 => b"00000_0000_00_000000000000", -- 0
 836 => b"00110_0000_01_000000000000", -- beq
 837 => b"00000_0000_00_001101110000", -- P2PLACEBOMB3
 838 => b"00000_0000_00_010001001101", -- load, gr0, P2BOMBCOUNT
 839 => b"00010_0000_01_000000000000", -- add, gr0
 840 => b"00000_0000_00_000000000001", -- 1
 841 => b"00001_0000_10_010001001101", -- store, gr0, P2BOMBCOUNT
 842 => b"00100_0000_01_000000000000", -- jump
 843 => b"00000_0000_00_001011000000", -- BTN2_R
 844 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 845 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 846 => b"00000_0011_00_010001010010", -- load, gr3, YPOS2
 847 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 848 => b"01000_0011_01_000000000000", -- mul, gr3
 849 => b"00000_0000_00_000000001111", -- 15
 850 => b"00010_0011_00_010001010001", -- add, gr3, XPOS2
 851 => b"10000_0011_00_000000000000", -- tpoint, gr3
 852 => b"01110_0010_00_000000000000", -- twrite, gr2
 853 => b"00000_0000_01_000000000000", -- load, gr0
 854 => b"00000_0000_00_000000000001", -- 1
 855 => b"00001_0000_10_010000111100", -- store, gr0, P2BOMB1ACTIVE
 856 => b"00001_0011_10_010000111010", -- store, gr3, P2BOMB1POS
 857 => b"00000_0000_01_000000000000", -- load, gr0
 858 => b"00000_0000_00_000000010000", -- 16
 859 => b"00001_0000_10_010000111011", -- store, gr0, P2BOMB1TIME
 860 => b"00100_0000_01_000000000000", -- jump
 861 => b"00000_0000_00_001101000110", -- P2INCREASEBOMBCOUNTER
 862 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 863 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 864 => b"00000_0011_00_010001010010", -- load, gr3, YPOS2
 865 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 866 => b"01000_0011_01_000000000000", -- mul, gr3
 867 => b"00000_0000_00_000000001111", -- 15
 868 => b"00010_0011_00_010001010001", -- add, gr3, XPOS2
 869 => b"10000_0011_00_000000000000", -- tpoint, gr3
 870 => b"01110_0010_00_000000000000", -- twrite, gr2
 871 => b"00000_0000_01_000000000000", -- load, gr0
 872 => b"00000_0000_00_000000000001", -- 1
 873 => b"00001_0000_10_010001000010", -- store, gr0, P2BOMB2ACTIVE
 874 => b"00001_0011_10_010001000000", -- store, gr3, P2BOMB2POS
 875 => b"00000_0000_01_000000000000", -- load, gr0
 876 => b"00000_0000_00_000000010000", -- 16
 877 => b"00001_0000_10_010001000001", -- store, gr0, P2BOMB2TIME
 878 => b"00100_0000_01_000000000000", -- jump
 879 => b"00000_0000_00_001101000110", -- P2INCREASEBOMBCOUNTER
 880 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 881 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 882 => b"00000_0011_00_010001010010", -- load, gr3, YPOS2
 883 => b"00000_0010_00_010001011010", -- load, gr2, EGG
 884 => b"01000_0011_01_000000000000", -- mul, gr3
 885 => b"00000_0000_00_000000001111", -- 15
 886 => b"00010_0011_00_010001010001", -- add, gr3, XPOS2
 887 => b"10000_0011_00_000000000000", -- tpoint, gr3
 888 => b"01110_0010_00_000000000000", -- twrite, gr2
 889 => b"00000_0000_01_000000000000", -- load, gr0
 890 => b"00000_0000_00_000000000001", -- 1
 891 => b"00001_0000_10_010001001000", -- store, gr0, P2BOMB3ACTIVE
 892 => b"00001_0011_10_010001000110", -- store, gr3, P2BOMB3POS
 893 => b"00000_0000_01_000000000000", -- load, gr0
 894 => b"00000_0000_00_000000010000", -- 16
 895 => b"00001_0000_10_010001000111", -- store, gr0, P2BOMB3TIME
 896 => b"00100_0000_01_000000000000", -- jump
 897 => b"00000_0000_00_001101000110", -- P2INCREASEBOMBCOUNTER
 898 => b"00000_0000_00_010000100110", -- load, gr0, P1DEAD
 899 => b"00011_0000_01_000000000000", -- sub, gr0
 900 => b"00000_0000_00_000000000001", -- 1
 901 => b"00110_0000_01_000000000000", -- beq
 902 => b"00000_0000_00_001110001111", -- J2
 903 => b"10001_0000_01_000000000000", -- joy1r
 904 => b"00000_0000_00_001110011110", -- P1R
 905 => b"10011_0000_01_000000000000", -- joy1l
 906 => b"00000_0000_00_001111000000", -- P1L
 907 => b"10010_0000_01_000000000000", -- joy1u
 908 => b"00000_0000_00_001110101111", -- P1U
 909 => b"10100_0000_01_000000000000", -- joy1d
 910 => b"00000_0000_00_001111010001", -- P1D
 911 => b"00000_0000_00_010000100111", -- load, gr0, P2DEAD
 912 => b"00011_0000_01_000000000000", -- sub, gr0
 913 => b"00000_0000_00_000000000001", -- 1
 914 => b"00110_0000_01_000000000000", -- beq
 915 => b"00000_0000_00_000001100110", -- CONTROL_R
 916 => b"10110_0000_01_000000000000", -- joy2r
 917 => b"00000_0000_00_001111100010", -- P2R
 918 => b"11000_0000_01_000000000000", -- joy2l
 919 => b"00000_0000_00_010000000100", -- P2L
 920 => b"10111_0000_01_000000000000", -- joy2u
 921 => b"00000_0000_00_001111110011", -- P2U
 922 => b"11001_0000_01_000000000000", -- joy2d
 923 => b"00000_0000_00_010000010101", -- P2D
 924 => b"00100_0000_01_000000000000", -- jump
 925 => b"00000_0000_00_000001100110", -- CONTROL_R
 926 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 927 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 928 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 929 => b"01000_0000_01_000000000000", -- mul, gr0
 930 => b"00000_0000_00_000000001111", -- 15
 931 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 932 => b"00010_0000_01_000000000000", -- add, gr0
 933 => b"00000_0000_00_000000000001", -- 1
 934 => b"10000_0000_00_000000000000", -- tpoint, gr0
 935 => b"01111_0001_00_000000000000", -- tread, gr1
 936 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
 937 => b"00111_0000_01_000000000000", -- bne
 938 => b"00000_0000_00_001110001011", -- J1
 939 => b"00010_1100_01_000000000000", -- add, gr12
 940 => b"00000_0000_00_000000000001", -- 1
 941 => b"00100_0000_01_000000000000", -- jump
 942 => b"00000_0000_00_001110001011", -- J1
 943 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 944 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 945 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 946 => b"00011_0000_01_000000000000", -- sub, gr0
 947 => b"00000_0000_00_000000000001", -- 1
 948 => b"01000_0000_01_000000000000", -- mul, gr0
 949 => b"00000_0000_00_000000001111", -- 15
 950 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 951 => b"10000_0000_00_000000000000", -- tpoint, gr0
 952 => b"01111_0001_00_000000000000", -- tread, gr1
 953 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
 954 => b"00111_0000_01_000000000000", -- bne
 955 => b"00000_0000_00_001110001111", -- J2
 956 => b"00011_1101_01_000000000000", -- sub, gr13
 957 => b"00000_0000_00_000000000001", -- 1
 958 => b"00100_0000_01_000000000000", -- jump
 959 => b"00000_0000_00_001110001111", -- J2
 960 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 961 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 962 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 963 => b"01000_0000_01_000000000000", -- mul, gr0
 964 => b"00000_0000_00_000000001111", -- 15
 965 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 966 => b"00011_0000_01_000000000000", -- sub, gr0
 967 => b"00000_0000_00_000000000001", -- 1
 968 => b"10000_0000_00_000000000000", -- tpoint, gr0
 969 => b"01111_0001_00_000000000000", -- tread, gr1
 970 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
 971 => b"00111_0000_01_000000000000", -- bne
 972 => b"00000_0000_00_001110001011", -- J1
 973 => b"00011_1100_01_000000000000", -- sub, gr12
 974 => b"00000_0000_00_000000000001", -- 1
 975 => b"00100_0000_01_000000000000", -- jump
 976 => b"00000_0000_00_001110001011", -- J1
 977 => b"00001_1100_10_010001001111", -- store, gr12, XPOS1
 978 => b"00001_1101_10_010001010000", -- store, gr13, YPOS1
 979 => b"00000_0000_00_010001010000", -- load, gr0, YPOS1
 980 => b"00010_0000_01_000000000000", -- add, gr0
 981 => b"00000_0000_00_000000000001", -- 1
 982 => b"01000_0000_01_000000000000", -- mul, gr0
 983 => b"00000_0000_00_000000001111", -- 15
 984 => b"00010_0000_00_010001001111", -- add, gr0, XPOS1
 985 => b"10000_0000_00_000000000000", -- tpoint, gr0
 986 => b"01111_0001_00_000000000000", -- tread, gr1
 987 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
 988 => b"00111_0000_01_000000000000", -- bne
 989 => b"00000_0000_00_001110001111", -- J2
 990 => b"00010_1101_01_000000000000", -- add, gr13
 991 => b"00000_0000_00_000000000001", -- 1
 992 => b"00100_0000_01_000000000000", -- jump
 993 => b"00000_0000_00_001110001111", -- J2
 994 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
 995 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
 996 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
 997 => b"01000_0000_01_000000000000", -- mul, gr0
 998 => b"00000_0000_00_000000001111", -- 15
 999 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
1000 => b"00010_0000_01_000000000000", -- add, gr0
1001 => b"00000_0000_00_000000000001", -- 1
1002 => b"10000_0000_00_000000000000", -- tpoint, gr0
1003 => b"01111_0001_00_000000000000", -- tread, gr1
1004 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
1005 => b"00111_0000_01_000000000000", -- bne
1006 => b"00000_0000_00_001110011000", -- J3
1007 => b"00010_1110_01_000000000000", -- add, gr14
1008 => b"00000_0000_00_000000000001", -- 1
1009 => b"00100_0000_01_000000000000", -- jump
1010 => b"00000_0000_00_001110011000", -- J3
1011 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
1012 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
1013 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
1014 => b"00011_0000_01_000000000000", -- sub, gr0
1015 => b"00000_0000_00_000000000001", -- 1
1016 => b"01000_0000_01_000000000000", -- mul, gr0
1017 => b"00000_0000_00_000000001111", -- 15
1018 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
1019 => b"10000_0000_00_000000000000", -- tpoint, gr0
1020 => b"01111_0001_00_000000000000", -- tread, gr1
1021 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
1022 => b"00111_0000_01_000000000000", -- bne
1023 => b"00000_0000_00_000001100110", -- CONTROL_R
1024 => b"00011_1111_01_000000000000", -- sub, gr15
1025 => b"00000_0000_00_000000000001", -- 1
1026 => b"00100_0000_01_000000000000", -- jump
1027 => b"00000_0000_00_000001100110", -- CONTROL_R
1028 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
1029 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
1030 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
1031 => b"01000_0000_01_000000000000", -- mul, gr0
1032 => b"00000_0000_00_000000001111", -- 15
1033 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
1034 => b"00011_0000_01_000000000000", -- sub, gr0
1035 => b"00000_0000_00_000000000001", -- 1
1036 => b"10000_0000_00_000000000000", -- tpoint, gr0
1037 => b"01111_0001_00_000000000000", -- tread, gr1
1038 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
1039 => b"00111_0000_01_000000000000", -- bne
1040 => b"00000_0000_00_001110011000", -- J3
1041 => b"00011_1110_01_000000000000", -- sub, gr14
1042 => b"00000_0000_00_000000000001", -- 1
1043 => b"00100_0000_01_000000000000", -- jump
1044 => b"00000_0000_00_001110011000", -- J3
1045 => b"00001_1110_10_010001010001", -- store, gr14, XPOS2
1046 => b"00001_1111_10_010001010010", -- store, gr15, YPOS2
1047 => b"00000_0000_00_010001010010", -- load, gr0, YPOS2
1048 => b"00010_0000_01_000000000000", -- add, gr0
1049 => b"00000_0000_00_000000000001", -- 1
1050 => b"01000_0000_01_000000000000", -- mul, gr0
1051 => b"00000_0000_00_000000001111", -- 15
1052 => b"00010_0000_00_010001010001", -- add, gr0, XPOS2
1053 => b"10000_0000_00_000000000000", -- tpoint, gr0
1054 => b"01111_0001_00_000000000000", -- tread, gr1
1055 => b"00011_0001_00_010001010110", -- sub, gr1, GRASS
1056 => b"00111_0000_01_000000000000", -- bne
1057 => b"00000_0000_00_000001100110", -- CONTROL_R
1058 => b"00010_1111_01_000000000000", -- add, gr15
1059 => b"00000_0000_00_000000000001", -- 1
1060 => b"00100_0000_01_000000000000", -- jump
1061 => b"00000_0000_00_000001100110", -- CONTROL_R
1062 => b"00000_0000_00_000000000000", -- 0
1063 => b"00000_0000_00_000000000000", -- 0
1064 => b"00000_0000_00_000000000000", -- 0
1065 => b"00000_0000_00_000000000000", -- 0
1066 => b"00000_0000_00_000000000000", -- 0
1067 => b"00000_0000_00_000000000000", -- 0
1068 => b"00000_0000_00_000000000000", -- 0
1069 => b"00000_0000_00_000000000000", -- 0
1070 => b"00000_0000_00_000000000000", -- 0
1071 => b"00000_0000_00_000000000000", -- 0
1072 => b"00000_0000_00_000000000000", -- 0
1073 => b"00000_0000_00_000000000000", -- 0
1074 => b"00000_0000_00_000000000000", -- 0
1075 => b"00000_0000_00_000000000000", -- 0
1076 => b"00000_0000_00_000000000000", -- 0
1077 => b"00000_0000_00_000000000000", -- 0
1078 => b"00000_0000_00_000000000000", -- 0
1079 => b"00000_0000_00_000000000000", -- 0
1080 => b"00000_0000_00_000000000000", -- 0
1081 => b"00000_0000_00_000000000000", -- 0
1082 => b"00000_0000_00_000000000000", -- 0
1083 => b"00000_0000_00_000000000000", -- 0
1084 => b"00000_0000_00_000000000000", -- 0
1085 => b"00000_0000_00_000000000000", -- 0
1086 => b"00000_0000_00_000000000000", -- 0
1087 => b"00000_0000_00_000000000000", -- 0
1088 => b"00000_0000_00_000000000000", -- 0
1089 => b"00000_0000_00_000000000000", -- 0
1090 => b"00000_0000_00_000000000000", -- 0
1091 => b"00000_0000_00_000000000000", -- 0
1092 => b"00000_0000_00_000000000000", -- 0
1093 => b"00000_0000_00_000000000000", -- 0
1094 => b"00000_0000_00_000000000000", -- 0
1095 => b"00000_0000_00_000000000000", -- 0
1096 => b"00000_0000_00_000000000000", -- 0
1097 => b"00000_0000_00_000000000000", -- 0
1098 => b"00000_0000_00_000000000000", -- 0
1099 => b"00000_0000_00_000000000000", -- 0
1100 => b"00000_0000_00_000000000000", -- 0
1101 => b"00000_0000_00_000000000000", -- 0
1102 => b"00000_0000_00_000000000011", -- 3
1103 => b"00000_0000_00_000000000000", -- 0
1104 => b"00000_0000_00_000000000000", -- 0
1105 => b"00000_0000_00_000000000000", -- 0
1106 => b"00000_0000_00_000000000000", -- 0
1107 => b"00000_0000_00_000000000000", -- 0
1108 => b"00000_0000_00_000000000000", -- 0
1109 => b"00000_0000_00_000000000000", -- 0
1110 => b"00000_0000_00_000000000000", -- 0
1111 => b"00000_0000_00_000000000001", -- 1
1112 => b"00000_0000_00_000000000010", -- 2
1113 => b"00000_0000_00_000000000011", -- 3
1114 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
