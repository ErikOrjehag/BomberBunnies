library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_0000_01_000000000000", -- load, gr0
   1 => b"00000_0000_00_000000000000", -- 0
   2 => b"00001_0000_10_010000001010", -- store, gr0, P1DEAD
   3 => b"00001_0000_10_010000001011", -- store, gr0, P2DEAD
   4 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMBCOUNT
   5 => b"00001_0000_10_010000110001", -- store, gr0, P2BOMBCOUNT
   6 => b"00000_1100_01_000000000000", -- load, gr12
   7 => b"00000_0000_00_000000000001", -- 1
   8 => b"00000_1101_01_000000000000", -- load, gr13
   9 => b"00000_0000_00_000000000001", -- 1
  10 => b"00000_1110_01_000000000000", -- load, gr14
  11 => b"00000_0000_00_000000001101", -- 13
  12 => b"00000_1111_01_000000000000", -- load, gr15
  13 => b"00000_0000_00_000000001011", -- 11
  14 => b"00001_0000_10_010000001100", -- store, gr0, P1BOMB1POS
  15 => b"00001_0000_10_010000001110", -- store, gr0, P1BOMB1ACTIVE
  16 => b"00001_0000_10_010000001101", -- store, gr0, P1BOMB1TIME
  17 => b"00001_0000_10_010000010010", -- store, gr0, P1BOMB2POS
  18 => b"00001_0000_10_010000010100", -- store, gr0, P1BOMB2ACTIVE
  19 => b"00001_0000_10_010000010011", -- store, gr0, P1BOMB2TIME
  20 => b"00001_0000_10_010000011000", -- store, gr0, P1BOMB3POS
  21 => b"00001_0000_10_010000011010", -- store, gr0, P1BOMB3ACTIVE
  22 => b"00001_0000_10_010000011001", -- store, gr0, P1BOMB3TIME
  23 => b"00001_0000_10_010000011110", -- store, gr0, P2BOMB1POS
  24 => b"00001_0000_10_010000100000", -- store, gr0, P2BOMB1ACTIVE
  25 => b"00001_0000_10_010000011111", -- store, gr0, P2BOMB1TIME
  26 => b"00001_0000_10_010000100100", -- store, gr0, P2BOMB2POS
  27 => b"00001_0000_10_010000100110", -- store, gr0, P2BOMB2ACTIVE
  28 => b"00001_0000_10_010000100101", -- store, gr0, P2BOMB2TIME
  29 => b"00001_0000_10_010000101010", -- store, gr0, P2BOMB3POS
  30 => b"00001_0000_10_010000101100", -- store, gr0, P2BOMB3ACTIVE
  31 => b"00001_0000_10_010000101011", -- store, gr0, P2BOMB3TIME
  32 => b"00001_0000_10_010000010001", -- store, gr0, P1EXPLOSION1POS
  33 => b"00001_0000_10_010000010000", -- store, gr0, P1EXPLOSION1ACTIVE
  34 => b"00001_0000_10_010000001111", -- store, gr0, P1EXPLOSION1TIME
  35 => b"00001_0000_10_010000010111", -- store, gr0, P1EXPLOSION2POS
  36 => b"00001_0000_10_010000010110", -- store, gr0, P1EXPLOSION2ACTIVE
  37 => b"00001_0000_10_010000010101", -- store, gr0, P1EXPLOSION2TIME
  38 => b"00001_0000_10_010000011101", -- store, gr0, P1EXPLOSION3POS
  39 => b"00001_0000_10_010000011100", -- store, gr0, P1EXPLOSION3ACTIVE
  40 => b"00001_0000_10_010000011011", -- store, gr0, P1EXPLOSION3TIME
  41 => b"00001_0000_10_010000100011", -- store, gr0, P2EXPLOSION1POS
  42 => b"00001_0000_10_010000100010", -- store, gr0, P2EXPLOSION1ACTIVE
  43 => b"00001_0000_10_010000100001", -- store, gr0, P2EXPLOSION1TIME
  44 => b"00001_0000_10_010000101001", -- store, gr0, P2EXPLOSION2POS
  45 => b"00001_0000_10_010000101000", -- store, gr0, P2EXPLOSION2ACTIVE
  46 => b"00001_0000_10_010000100111", -- store, gr0, P2EXPLOSION2TIME
  47 => b"00001_0000_10_010000101111", -- store, gr0, P2EXPLOSION3POS
  48 => b"00001_0000_10_010000101110", -- store, gr0, P2EXPLOSION3ACTIVE
  49 => b"00001_0000_10_010000101101", -- store, gr0, P2EXPLOSION3TIME
  50 => b"00000_0000_01_000000000000", -- load, gr0
  51 => b"00000_0000_00_000000000000", -- 0
  52 => b"00000_0011_01_000000000000", -- load, gr3
  53 => b"00000_0000_00_000011000011", -- 195
  54 => b"00001_0000_10_010000110111", -- store, gr0, MOVE
  55 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
  56 => b"00001_0011_10_010000110111", -- store, gr3, MOVE
  57 => b"00011_0010_00_010000110111", -- sub, gr2, MOVE
  58 => b"00110_0000_01_000000000000", -- beq
  59 => b"00000_0000_00_000001000111", -- INITEND
  60 => b"10000_0000_00_000000000000", -- tpoint, gr0
  61 => b"01111_0001_00_000000000000", -- tread, gr1
  62 => b"00011_0001_00_010000111011", -- sub, gr1, WALL
  63 => b"00110_0000_01_000000000000", -- beq
  64 => b"00000_0000_00_000001000011", -- INCREASE
  65 => b"00000_0001_00_010000111100", -- load, gr1, BREAKABLE
  66 => b"01110_0001_00_000000000000", -- twrite, gr1
  67 => b"00010_0000_01_000000000000", -- add, gr0
  68 => b"00000_0000_00_000000000001", -- 1
  69 => b"00100_0000_01_000000000000", -- jump
  70 => b"00000_0000_00_000000110110", -- INITLOOP
  71 => b"00000_0000_00_010000111010", -- load, gr0, GRASS
  72 => b"00000_0001_01_000000000000", -- load, gr1
  73 => b"00000_0000_00_000000010000", -- 16
  74 => b"10000_0001_00_000000000000", -- tpoint, gr1
  75 => b"01110_0000_00_000000000000", -- twrite, gr0
  76 => b"00010_0001_01_000000000000", -- add, gr1
  77 => b"00000_0000_00_000000000001", -- 1
  78 => b"10000_0001_00_000000000000", -- tpoint, gr1
  79 => b"01110_0000_00_000000000000", -- twrite, gr0
  80 => b"00010_0001_01_000000000000", -- add, gr1
  81 => b"00000_0000_00_000000001110", -- 14
  82 => b"10000_0001_00_000000000000", -- tpoint, gr1
  83 => b"01110_0000_00_000000000000", -- twrite, gr0
  84 => b"00000_0001_01_000000000000", -- load, gr1
  85 => b"00000_0000_00_000010110010", -- 178
  86 => b"10000_0001_00_000000000000", -- tpoint, gr1
  87 => b"01110_0000_00_000000000000", -- twrite, gr0
  88 => b"00011_0001_01_000000000000", -- sub, gr1
  89 => b"00000_0000_00_000000000001", -- 1
  90 => b"10000_0001_00_000000000000", -- tpoint, gr1
  91 => b"01110_0000_00_000000000000", -- twrite, gr0
  92 => b"00011_0001_01_000000000000", -- sub, gr1
  93 => b"00000_0000_00_000000001110", -- 14
  94 => b"10000_0001_00_000000000000", -- tpoint, gr1
  95 => b"01110_0000_00_000000000000", -- twrite, gr0
  96 => b"00100_0000_01_000000000000", -- jump
  97 => b"00000_0000_00_000010101000", -- CHECKDEATH
  98 => b"00100_0000_01_000000000000", -- jump
  99 => b"00000_0000_00_000001101110", -- CHECKBOMBDEATH
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_001101100110", -- CONTROL
 102 => b"00100_0000_01_000000000000", -- jump
 103 => b"00000_0000_00_001010100000", -- BUTTON
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000110010001", -- TICKBOMBS
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000011001010", -- TICKEXPLOSIONS
 108 => b"00100_0000_01_000000000000", -- jump
 109 => b"00000_0000_00_000001100000", -- MAIN
 110 => b"00000_0010_01_000000000000", -- load, gr2
 111 => b"00000_0000_00_000000000001", -- 1
 112 => b"00000_0000_00_010000001100", -- load, gr0, P1BOMB1POS
 113 => b"10000_0000_00_000000000000", -- tpoint, gr0
 114 => b"01111_0001_00_000000000000", -- tread, gr1
 115 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 116 => b"00110_0000_01_000000000000", -- beq
 117 => b"00000_0000_00_000010010110", -- P1BOMB1DETONATE
 118 => b"00000_0000_00_010000010010", -- load, gr0, P1BOMB2POS
 119 => b"10000_0000_00_000000000000", -- tpoint, gr0
 120 => b"01111_0001_00_000000000000", -- tread, gr1
 121 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 122 => b"00110_0000_01_000000000000", -- beq
 123 => b"00000_0000_00_000010011001", -- P1BOMB2DETONATE
 124 => b"00000_0000_00_010000011000", -- load, gr0, P1BOMB3POS
 125 => b"10000_0000_00_000000000000", -- tpoint, gr0
 126 => b"01111_0001_00_000000000000", -- tread, gr1
 127 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 128 => b"00110_0000_01_000000000000", -- beq
 129 => b"00000_0000_00_000010011100", -- P1BOMB3DETONATE
 130 => b"00000_0000_00_010000011110", -- load, gr0, P2BOMB1POS
 131 => b"10000_0000_00_000000000000", -- tpoint, gr0
 132 => b"01111_0001_00_000000000000", -- tread, gr1
 133 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 134 => b"00110_0000_01_000000000000", -- beq
 135 => b"00000_0000_00_000010011111", -- P2BOMB1DETONATE
 136 => b"00000_0000_00_010000100100", -- load, gr0, P2BOMB2POS
 137 => b"10000_0000_00_000000000000", -- tpoint, gr0
 138 => b"01111_0001_00_000000000000", -- tread, gr1
 139 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 140 => b"00110_0000_01_000000000000", -- beq
 141 => b"00000_0000_00_000010100010", -- P2BOMB2DETONATE
 142 => b"00000_0000_00_010000101010", -- load, gr0, P2BOMB3POS
 143 => b"10000_0000_00_000000000000", -- tpoint, gr0
 144 => b"01111_0001_00_000000000000", -- tread, gr1
 145 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 146 => b"00110_0000_01_000000000000", -- beq
 147 => b"00000_0000_00_000010100101", -- P2BOMB3DETONATE
 148 => b"00100_0000_01_000000000000", -- jump
 149 => b"00000_0000_00_000001100100", -- CHECKBOMBDEATH_R
 150 => b"00001_0010_10_010000001101", -- store, gr2, P1BOMB1TIME
 151 => b"00100_0000_01_000000000000", -- jump
 152 => b"00000_0000_00_000001110110", -- P1BOMB1DETONATE_R
 153 => b"00001_0010_10_010000010011", -- store, gr2, P1BOMB2TIME
 154 => b"00100_0000_01_000000000000", -- jump
 155 => b"00000_0000_00_000001111100", -- P1BOMB2DETONATE_R
 156 => b"00001_0010_10_010000011001", -- store, gr2, P1BOMB3TIME
 157 => b"00100_0000_01_000000000000", -- jump
 158 => b"00000_0000_00_000010000010", -- P1BOMB3DETONATE_R
 159 => b"00001_0010_10_010000011111", -- store, gr2, P2BOMB1TIME
 160 => b"00100_0000_01_000000000000", -- jump
 161 => b"00000_0000_00_000010001000", -- P2BOMB1DETONATE_R
 162 => b"00001_0010_10_010000100101", -- store, gr2, P2BOMB2TIME
 163 => b"00100_0000_01_000000000000", -- jump
 164 => b"00000_0000_00_000010001110", -- P2BOMB2DETONATE_R
 165 => b"00001_0010_10_010000101011", -- store, gr2, P2BOMB3TIME
 166 => b"00100_0000_01_000000000000", -- jump
 167 => b"00000_0000_00_000010010100", -- P2BOMB3DETONATE_R
 168 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 169 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 170 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 171 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 172 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 173 => b"01000_0000_01_000000000000", -- mul, gr0
 174 => b"00000_0000_00_000000001111", -- 15
 175 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 176 => b"10000_0000_00_000000000000", -- tpoint, gr0
 177 => b"01111_0001_00_000000000000", -- tread, gr1
 178 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 179 => b"00110_0000_01_000000000000", -- beq
 180 => b"00000_0000_00_000011000000", -- P1DEATH
 181 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
 182 => b"01000_0000_01_000000000000", -- mul, gr0
 183 => b"00000_0000_00_000000001111", -- 15
 184 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
 185 => b"10000_0000_00_000000000000", -- tpoint, gr0
 186 => b"01111_0001_00_000000000000", -- tread, gr1
 187 => b"00011_0001_00_010000111101", -- sub, gr1, EXPLOSION
 188 => b"00110_0000_01_000000000000", -- beq
 189 => b"00000_0000_00_000011000101", -- P2DEATH
 190 => b"00100_0000_01_000000000000", -- jump
 191 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 192 => b"00000_0000_01_000000000000", -- load, gr0
 193 => b"00000_0000_00_000000000001", -- 1
 194 => b"00001_0000_10_010000001010", -- store, gr0, P1DEAD
 195 => b"00100_0000_01_000000000000", -- jump
 196 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 197 => b"00000_0000_01_000000000000", -- load, gr0
 198 => b"00000_0000_00_000000000001", -- 1
 199 => b"00001_0000_10_010000001011", -- store, gr0, P2DEAD
 200 => b"00100_0000_01_000000000000", -- jump
 201 => b"00000_0000_00_000001100010", -- CHECKDEATH_R
 202 => b"00000_0000_00_010000010000", -- load, gr0, P1EXPLOSION1ACTIVE
 203 => b"00011_0000_01_000000000000", -- sub, gr0
 204 => b"00000_0000_00_000000000001", -- 1
 205 => b"00111_0000_01_000000000000", -- bne
 206 => b"00000_0000_00_000011011000", -- P1EXPLOSION2
 207 => b"00000_0000_00_010000001111", -- load, gr0, P1EXPLOSION1TIME
 208 => b"00011_0000_01_000000000000", -- sub, gr0
 209 => b"00000_0000_00_000000000001", -- 1
 210 => b"00001_0000_10_010000001111", -- store, gr0, P1EXPLOSION1TIME
 211 => b"00000_0000_01_000000000000", -- load, gr0
 212 => b"00000_0000_00_000000000000", -- 0
 213 => b"00011_0000_00_010000001111", -- sub, gr0, P1EXPLOSION1TIME
 214 => b"00110_0000_01_000000000000", -- beq
 215 => b"00000_0000_00_000100100000", -- P1EXPLOSION1FADE
 216 => b"00000_0000_00_010000010110", -- load, gr0, P1EXPLOSION2ACTIVE
 217 => b"00011_0000_01_000000000000", -- sub, gr0
 218 => b"00000_0000_00_000000000001", -- 1
 219 => b"00111_0000_01_000000000000", -- bne
 220 => b"00000_0000_00_000011100110", -- P1EXPLOSION3
 221 => b"00000_0000_00_010000010101", -- load, gr0, P1EXPLOSION2TIME
 222 => b"00011_0000_01_000000000000", -- sub, gr0
 223 => b"00000_0000_00_000000000001", -- 1
 224 => b"00001_0000_10_010000010101", -- store, gr0, P1EXPLOSION2TIME
 225 => b"00000_0000_01_000000000000", -- load, gr0
 226 => b"00000_0000_00_000000000000", -- 0
 227 => b"00011_0000_00_010000010101", -- sub, gr0, P1EXPLOSION2TIME
 228 => b"00110_0000_01_000000000000", -- beq
 229 => b"00000_0000_00_000100100110", -- P1EXPLOSION2FADE
 230 => b"00000_0000_00_010000011100", -- load, gr0, P1EXPLOSION3ACTIVE
 231 => b"00011_0000_01_000000000000", -- sub, gr0
 232 => b"00000_0000_00_000000000001", -- 1
 233 => b"00111_0000_01_000000000000", -- bne
 234 => b"00000_0000_00_000011110100", -- P2EXPLOSION1
 235 => b"00000_0000_00_010000011011", -- load, gr0, P1EXPLOSION3TIME
 236 => b"00011_0000_01_000000000000", -- sub, gr0
 237 => b"00000_0000_00_000000000001", -- 1
 238 => b"00001_0000_10_010000011011", -- store, gr0, P1EXPLOSION3TIME
 239 => b"00000_0000_01_000000000000", -- load, gr0
 240 => b"00000_0000_00_000000000000", -- 0
 241 => b"00011_0000_00_010000011011", -- sub, gr0, P1EXPLOSION3TIME
 242 => b"00110_0000_01_000000000000", -- beq
 243 => b"00000_0000_00_000100101100", -- P1EXPLOSION3FADE
 244 => b"00000_0000_00_010000100010", -- load, gr0, P2EXPLOSION1ACTIVE
 245 => b"00011_0000_01_000000000000", -- sub, gr0
 246 => b"00000_0000_00_000000000001", -- 1
 247 => b"00111_0000_01_000000000000", -- bne
 248 => b"00000_0000_00_000100000010", -- P2EXPLOSION2
 249 => b"00000_0000_00_010000100001", -- load, gr0, P2EXPLOSION1TIME
 250 => b"00011_0000_01_000000000000", -- sub, gr0
 251 => b"00000_0000_00_000000000001", -- 1
 252 => b"00001_0000_10_010000100001", -- store, gr0, P2EXPLOSION1TIME
 253 => b"00000_0000_01_000000000000", -- load, gr0
 254 => b"00000_0000_00_000000000000", -- 0
 255 => b"00011_0000_00_010000100001", -- sub, gr0, P2EXPLOSION1TIME
 256 => b"00110_0000_01_000000000000", -- beq
 257 => b"00000_0000_00_000100110010", -- P2EXPLOSION1FADE
 258 => b"00000_0000_00_010000101000", -- load, gr0, P2EXPLOSION2ACTIVE
 259 => b"00011_0000_01_000000000000", -- sub, gr0
 260 => b"00000_0000_00_000000000001", -- 1
 261 => b"00111_0000_01_000000000000", -- bne
 262 => b"00000_0000_00_000100010000", -- P2EXPLOSION3
 263 => b"00000_0000_00_010000100111", -- load, gr0, P2EXPLOSION2TIME
 264 => b"00011_0000_01_000000000000", -- sub, gr0
 265 => b"00000_0000_00_000000000001", -- 1
 266 => b"00001_0000_10_010000100111", -- store, gr0, P2EXPLOSION2TIME
 267 => b"00000_0000_01_000000000000", -- load, gr0
 268 => b"00000_0000_00_000000000000", -- 0
 269 => b"00011_0000_00_010000100111", -- sub, gr0, P2EXPLOSION2TIME
 270 => b"00110_0000_01_000000000000", -- beq
 271 => b"00000_0000_00_000100111000", -- P2EXPLOSION2FADE
 272 => b"00000_0000_00_010000101110", -- load, gr0, P2EXPLOSION3ACTIVE
 273 => b"00011_0000_01_000000000000", -- sub, gr0
 274 => b"00000_0000_00_000000000001", -- 1
 275 => b"00111_0000_01_000000000000", -- bne
 276 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 277 => b"00000_0000_00_010000101101", -- load, gr0, P2EXPLOSION3TIME
 278 => b"00011_0000_01_000000000000", -- sub, gr0
 279 => b"00000_0000_00_000000000001", -- 1
 280 => b"00001_0000_10_010000101101", -- store, gr0, P2EXPLOSION3TIME
 281 => b"00000_0000_01_000000000000", -- load, gr0
 282 => b"00000_0000_00_000000000000", -- 0
 283 => b"00011_0000_00_010000101101", -- sub, gr0, P2EXPLOSION3TIME
 284 => b"00110_0000_01_000000000000", -- beq
 285 => b"00000_0000_00_000100111110", -- P2EXPLOSION3FADE
 286 => b"00100_0000_01_000000000000", -- jump
 287 => b"00000_0000_00_000001101100", -- TICKEXPLOSIONS_R
 288 => b"00000_0000_01_000000000000", -- load, gr0
 289 => b"00000_0000_00_000000000000", -- 0
 290 => b"00001_0000_10_010000010000", -- store, gr0, P1EXPLOSION1ACTIVE
 291 => b"00000_0100_00_010000010001", -- load, gr4, P1EXPLOSION1POS
 292 => b"00100_0000_01_000000000000", -- jump
 293 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 294 => b"00000_0000_01_000000000000", -- load, gr0
 295 => b"00000_0000_00_000000000000", -- 0
 296 => b"00001_0000_10_010000010110", -- store, gr0, P1EXPLOSION2ACTIVE
 297 => b"00000_0100_00_010000010111", -- load, gr4, P1EXPLOSION2POS
 298 => b"00100_0000_01_000000000000", -- jump
 299 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 300 => b"00000_0000_01_000000000000", -- load, gr0
 301 => b"00000_0000_00_000000000000", -- 0
 302 => b"00001_0000_10_010000011100", -- store, gr0, P1EXPLOSION3ACTIVE
 303 => b"00000_0100_00_010000011101", -- load, gr4, P1EXPLOSION3POS
 304 => b"00100_0000_01_000000000000", -- jump
 305 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 306 => b"00000_0000_01_000000000000", -- load, gr0
 307 => b"00000_0000_00_000000000000", -- 0
 308 => b"00001_0000_10_010000100010", -- store, gr0, P2EXPLOSION1ACTIVE
 309 => b"00000_0100_00_010000100011", -- load, gr4, P2EXPLOSION1POS
 310 => b"00100_0000_01_000000000000", -- jump
 311 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 312 => b"00000_0000_01_000000000000", -- load, gr0
 313 => b"00000_0000_00_000000000000", -- 0
 314 => b"00001_0000_10_010000101000", -- store, gr0, P2EXPLOSION2ACTIVE
 315 => b"00000_0100_00_010000101001", -- load, gr4, P2EXPLOSION2POS
 316 => b"00100_0000_01_000000000000", -- jump
 317 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 318 => b"00000_0000_01_000000000000", -- load, gr0
 319 => b"00000_0000_00_000000000000", -- 0
 320 => b"00001_0000_10_010000101110", -- store, gr0, P2EXPLOSION3ACTIVE
 321 => b"00000_0100_00_010000101111", -- load, gr4, P2EXPLOSION3POS
 322 => b"00100_0000_01_000000000000", -- jump
 323 => b"00000_0000_00_000101000100", -- FADEEXPLOSION
 324 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 325 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 326 => b"00000_0011_00_010000111010", -- load, gr3, GRASS
 327 => b"10000_0010_00_000000000000", -- tpoint, gr2
 328 => b"01110_0011_00_000000000000", -- twrite, gr3
 329 => b"00010_0010_01_000000000000", -- add, gr2
 330 => b"00000_0000_00_000000000001", -- 1
 331 => b"10000_0010_00_000000000000", -- tpoint, gr2
 332 => b"01111_0000_00_000000000000", -- tread, gr0
 333 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 334 => b"00111_0000_01_000000000000", -- bne
 335 => b"00000_0000_00_000101011001", -- FADELEFT
 336 => b"01110_0011_00_000000000000", -- twrite, gr3
 337 => b"00010_0010_01_000000000000", -- add, gr2
 338 => b"00000_0000_00_000000000001", -- 1
 339 => b"10000_0010_00_000000000000", -- tpoint, gr2
 340 => b"01111_0000_00_000000000000", -- tread, gr0
 341 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 342 => b"00111_0000_01_000000000000", -- bne
 343 => b"00000_0000_00_000101011001", -- FADELEFT
 344 => b"01110_0011_00_000000000000", -- twrite, gr3
 345 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 346 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 347 => b"00011_0010_01_000000000000", -- sub, gr2
 348 => b"00000_0000_00_000000000001", -- 1
 349 => b"10000_0010_00_000000000000", -- tpoint, gr2
 350 => b"01111_0000_00_000000000000", -- tread, gr0
 351 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 352 => b"00111_0000_01_000000000000", -- bne
 353 => b"00000_0000_00_000101101011", -- FADEDOWN
 354 => b"01110_0011_00_000000000000", -- twrite, gr3
 355 => b"00011_0010_01_000000000000", -- sub, gr2
 356 => b"00000_0000_00_000000000001", -- 1
 357 => b"10000_0010_00_000000000000", -- tpoint, gr2
 358 => b"01111_0000_00_000000000000", -- tread, gr0
 359 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 360 => b"00111_0000_01_000000000000", -- bne
 361 => b"00000_0000_00_000101101011", -- FADEDOWN
 362 => b"01110_0011_00_000000000000", -- twrite, gr3
 363 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 364 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 365 => b"00010_0010_01_000000000000", -- add, gr2
 366 => b"00000_0000_00_000000001111", -- 15
 367 => b"10000_0010_00_000000000000", -- tpoint, gr2
 368 => b"01111_0000_00_000000000000", -- tread, gr0
 369 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 370 => b"00111_0000_01_000000000000", -- bne
 371 => b"00000_0000_00_000101111101", -- FADEUP
 372 => b"01110_0011_00_000000000000", -- twrite, gr3
 373 => b"00010_0010_01_000000000000", -- add, gr2
 374 => b"00000_0000_00_000000001111", -- 15
 375 => b"10000_0010_00_000000000000", -- tpoint, gr2
 376 => b"01111_0000_00_000000000000", -- tread, gr0
 377 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 378 => b"00111_0000_01_000000000000", -- bne
 379 => b"00000_0000_00_000101111101", -- FADEUP
 380 => b"01110_0011_00_000000000000", -- twrite, gr3
 381 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 382 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 383 => b"00011_0010_01_000000000000", -- sub, gr2
 384 => b"00000_0000_00_000000001111", -- 15
 385 => b"10000_0010_00_000000000000", -- tpoint, gr2
 386 => b"01111_0000_00_000000000000", -- tread, gr0
 387 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 388 => b"00111_0000_01_000000000000", -- bne
 389 => b"00000_0000_00_000011001010", -- TICKEXPLOSIONS
 390 => b"01110_0011_00_000000000000", -- twrite, gr3
 391 => b"00011_0010_01_000000000000", -- sub, gr2
 392 => b"00000_0000_00_000000001111", -- 15
 393 => b"10000_0010_00_000000000000", -- tpoint, gr2
 394 => b"01111_0000_00_000000000000", -- tread, gr0
 395 => b"00011_0000_00_010000111101", -- sub, gr0, EXPLOSION
 396 => b"00111_0000_01_000000000000", -- bne
 397 => b"00000_0000_00_000011001010", -- TICKEXPLOSIONS
 398 => b"01110_0011_00_000000000000", -- twrite, gr3
 399 => b"00100_0000_01_000000000000", -- jump
 400 => b"00000_0000_00_000011001010", -- TICKEXPLOSIONS
 401 => b"00000_0000_00_010000001110", -- load, gr0, P1BOMB1ACTIVE
 402 => b"00011_0000_01_000000000000", -- sub, gr0
 403 => b"00000_0000_00_000000000001", -- 1
 404 => b"00111_0000_01_000000000000", -- bne
 405 => b"00000_0000_00_000110011111", -- P1BOMB2
 406 => b"00000_0000_00_010000001101", -- load, gr0, P1BOMB1TIME
 407 => b"00011_0000_01_000000000000", -- sub, gr0
 408 => b"00000_0000_00_000000000001", -- 1
 409 => b"00001_0000_10_010000001101", -- store, gr0, P1BOMB1TIME
 410 => b"00000_0000_01_000000000000", -- load, gr0
 411 => b"00000_0000_00_000000000000", -- 0
 412 => b"00011_0000_00_010000001101", -- sub, gr0, P1BOMB1TIME
 413 => b"00110_0000_01_000000000000", -- beq
 414 => b"00000_0000_00_000111100111", -- P1EXPLOSION1INIT
 415 => b"00000_0000_00_010000010100", -- load, gr0, P1BOMB2ACTIVE
 416 => b"00011_0000_01_000000000000", -- sub, gr0
 417 => b"00000_0000_00_000000000001", -- 1
 418 => b"00111_0000_01_000000000000", -- bne
 419 => b"00000_0000_00_000110101101", -- P1BOMB3
 420 => b"00000_0000_00_010000010011", -- load, gr0, P1BOMB2TIME
 421 => b"00011_0000_01_000000000000", -- sub, gr0
 422 => b"00000_0000_00_000000000001", -- 1
 423 => b"00001_0000_10_010000010011", -- store, gr0, P1BOMB2TIME
 424 => b"00000_0000_01_000000000000", -- load, gr0
 425 => b"00000_0000_00_000000000000", -- 0
 426 => b"00011_0000_00_010000010011", -- sub, gr0, P1BOMB2TIME
 427 => b"00110_0000_01_000000000000", -- beq
 428 => b"00000_0000_00_000111111001", -- P1EXPLOSION2INIT
 429 => b"00000_0000_00_010000011010", -- load, gr0, P1BOMB3ACTIVE
 430 => b"00011_0000_01_000000000000", -- sub, gr0
 431 => b"00000_0000_00_000000000001", -- 1
 432 => b"00111_0000_01_000000000000", -- bne
 433 => b"00000_0000_00_000110111011", -- P2BOMB1
 434 => b"00000_0000_00_010000011001", -- load, gr0, P1BOMB3TIME
 435 => b"00011_0000_01_000000000000", -- sub, gr0
 436 => b"00000_0000_00_000000000001", -- 1
 437 => b"00001_0000_10_010000011001", -- store, gr0, P1BOMB3TIME
 438 => b"00000_0000_01_000000000000", -- load, gr0
 439 => b"00000_0000_00_000000000000", -- 0
 440 => b"00011_0000_00_010000011001", -- sub, gr0, P1BOMB3TIME
 441 => b"00110_0000_01_000000000000", -- beq
 442 => b"00000_0000_00_001000001011", -- P1EXPLOSION3INIT
 443 => b"00000_0000_00_010000100000", -- load, gr0, P2BOMB1ACTIVE
 444 => b"00011_0000_01_000000000000", -- sub, gr0
 445 => b"00000_0000_00_000000000001", -- 1
 446 => b"00111_0000_01_000000000000", -- bne
 447 => b"00000_0000_00_000111001001", -- P2BOMB2
 448 => b"00000_0000_00_010000011111", -- load, gr0, P2BOMB1TIME
 449 => b"00011_0000_01_000000000000", -- sub, gr0
 450 => b"00000_0000_00_000000000001", -- 1
 451 => b"00001_0000_10_010000011111", -- store, gr0, P2BOMB1TIME
 452 => b"00000_0000_01_000000000000", -- load, gr0
 453 => b"00000_0000_00_000000000000", -- 0
 454 => b"00011_0000_00_010000011111", -- sub, gr0, P2BOMB1TIME
 455 => b"00110_0000_01_000000000000", -- beq
 456 => b"00000_0000_00_001000011101", -- P2EXPLOSION1INIT
 457 => b"00000_0000_00_010000100110", -- load, gr0, P2BOMB2ACTIVE
 458 => b"00011_0000_01_000000000000", -- sub, gr0
 459 => b"00000_0000_00_000000000001", -- 1
 460 => b"00111_0000_01_000000000000", -- bne
 461 => b"00000_0000_00_000111010111", -- P2BOMB3
 462 => b"00000_0000_00_010000100101", -- load, gr0, P2BOMB2TIME
 463 => b"00011_0000_01_000000000000", -- sub, gr0
 464 => b"00000_0000_00_000000000001", -- 1
 465 => b"00001_0000_10_010000100101", -- store, gr0, P2BOMB2TIME
 466 => b"00000_0000_01_000000000000", -- load, gr0
 467 => b"00000_0000_00_000000000000", -- 0
 468 => b"00011_0000_00_010000100101", -- sub, gr0, P2BOMB2TIME
 469 => b"00110_0000_01_000000000000", -- beq
 470 => b"00000_0000_00_001000101111", -- P2EXPLOSION2INIT
 471 => b"00000_0000_00_010000101100", -- load, gr0, P2BOMB3ACTIVE
 472 => b"00011_0000_01_000000000000", -- sub, gr0
 473 => b"00000_0000_00_000000000001", -- 1
 474 => b"00111_0000_01_000000000000", -- bne
 475 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 476 => b"00000_0000_00_010000101011", -- load, gr0, P2BOMB3TIME
 477 => b"00011_0000_01_000000000000", -- sub, gr0
 478 => b"00000_0000_00_000000000001", -- 1
 479 => b"00001_0000_10_010000101011", -- store, gr0, P2BOMB3TIME
 480 => b"00000_0000_01_000000000000", -- load, gr0
 481 => b"00000_0000_00_000000000000", -- 0
 482 => b"00011_0000_00_010000101011", -- sub, gr0, P2BOMB3TIME
 483 => b"00110_0000_01_000000000000", -- beq
 484 => b"00000_0000_00_001001000001", -- P2EXPLOSION3INIT
 485 => b"00100_0000_01_000000000000", -- jump
 486 => b"00000_0000_00_000001101010", -- TICKBOMBS_R
 487 => b"00000_0000_01_000000000000", -- load, gr0
 488 => b"00000_0000_00_000000000000", -- 0
 489 => b"00001_0000_10_010000001110", -- store, gr0, P1BOMB1ACTIVE
 490 => b"00000_0000_00_010000001100", -- load, gr0, P1BOMB1POS
 491 => b"00001_0000_10_010000010001", -- store, gr0, P1EXPLOSION1POS
 492 => b"00000_0000_01_000000000000", -- load, gr0
 493 => b"00000_0000_00_000000000001", -- 1
 494 => b"00001_0000_10_010000010000", -- store, gr0, P1EXPLOSION1ACTIVE
 495 => b"00000_0000_01_000000000000", -- load, gr0
 496 => b"00000_0000_00_000000000010", -- 2
 497 => b"00001_0000_10_010000001111", -- store, gr0, P1EXPLOSION1TIME
 498 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMBCOUNT
 499 => b"00011_0000_01_000000000000", -- sub, gr0
 500 => b"00000_0000_00_000000000001", -- 1
 501 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMBCOUNT
 502 => b"00000_0100_00_010000001100", -- load, gr4, P1BOMB1POS
 503 => b"00100_0000_01_000000000000", -- jump
 504 => b"00000_0000_00_001001010011", -- EXPLODE
 505 => b"00000_0000_01_000000000000", -- load, gr0
 506 => b"00000_0000_00_000000000000", -- 0
 507 => b"00001_0000_10_010000010100", -- store, gr0, P1BOMB2ACTIVE
 508 => b"00000_0000_00_010000010010", -- load, gr0, P1BOMB2POS
 509 => b"00001_0000_10_010000010111", -- store, gr0, P1EXPLOSION2POS
 510 => b"00000_0000_01_000000000000", -- load, gr0
 511 => b"00000_0000_00_000000000001", -- 1
 512 => b"00001_0000_10_010000010110", -- store, gr0, P1EXPLOSION2ACTIVE
 513 => b"00000_0000_01_000000000000", -- load, gr0
 514 => b"00000_0000_00_000000000010", -- 2
 515 => b"00001_0000_10_010000010101", -- store, gr0, P1EXPLOSION2TIME
 516 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMBCOUNT
 517 => b"00011_0000_01_000000000000", -- sub, gr0
 518 => b"00000_0000_00_000000000001", -- 1
 519 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMBCOUNT
 520 => b"00000_0100_00_010000010010", -- load, gr4, P1BOMB2POS
 521 => b"00100_0000_01_000000000000", -- jump
 522 => b"00000_0000_00_001001010011", -- EXPLODE
 523 => b"00000_0000_01_000000000000", -- load, gr0
 524 => b"00000_0000_00_000000000000", -- 0
 525 => b"00001_0000_10_010000011010", -- store, gr0, P1BOMB3ACTIVE
 526 => b"00000_0000_00_010000011000", -- load, gr0, P1BOMB3POS
 527 => b"00001_0000_10_010000011101", -- store, gr0, P1EXPLOSION3POS
 528 => b"00000_0000_01_000000000000", -- load, gr0
 529 => b"00000_0000_00_000000000001", -- 1
 530 => b"00001_0000_10_010000011100", -- store, gr0, P1EXPLOSION3ACTIVE
 531 => b"00000_0000_01_000000000000", -- load, gr0
 532 => b"00000_0000_00_000000000010", -- 2
 533 => b"00001_0000_10_010000011011", -- store, gr0, P1EXPLOSION3TIME
 534 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMBCOUNT
 535 => b"00011_0000_01_000000000000", -- sub, gr0
 536 => b"00000_0000_00_000000000001", -- 1
 537 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMBCOUNT
 538 => b"00000_0100_00_010000011000", -- load, gr4, P1BOMB3POS
 539 => b"00100_0000_01_000000000000", -- jump
 540 => b"00000_0000_00_001001010011", -- EXPLODE
 541 => b"00000_0000_01_000000000000", -- load, gr0
 542 => b"00000_0000_00_000000000000", -- 0
 543 => b"00001_0000_10_010000100000", -- store, gr0, P2BOMB1ACTIVE
 544 => b"00000_0000_00_010000011110", -- load, gr0, P2BOMB1POS
 545 => b"00001_0000_10_010000100011", -- store, gr0, P2EXPLOSION1POS
 546 => b"00000_0000_01_000000000000", -- load, gr0
 547 => b"00000_0000_00_000000000001", -- 1
 548 => b"00001_0000_10_010000100010", -- store, gr0, P2EXPLOSION1ACTIVE
 549 => b"00000_0000_01_000000000000", -- load, gr0
 550 => b"00000_0000_00_000000000010", -- 2
 551 => b"00001_0000_10_010000100001", -- store, gr0, P2EXPLOSION1TIME
 552 => b"00000_0000_00_010000110001", -- load, gr0, P2BOMBCOUNT
 553 => b"00011_0000_01_000000000000", -- sub, gr0
 554 => b"00000_0000_00_000000000001", -- 1
 555 => b"00001_0000_10_010000110001", -- store, gr0, P2BOMBCOUNT
 556 => b"00000_0100_00_010000011110", -- load, gr4, P2BOMB1POS
 557 => b"00100_0000_01_000000000000", -- jump
 558 => b"00000_0000_00_001001010011", -- EXPLODE
 559 => b"00000_0000_01_000000000000", -- load, gr0
 560 => b"00000_0000_00_000000000000", -- 0
 561 => b"00001_0000_10_010000100110", -- store, gr0, P2BOMB2ACTIVE
 562 => b"00000_0000_00_010000100100", -- load, gr0, P2BOMB2POS
 563 => b"00001_0000_10_010000101001", -- store, gr0, P2EXPLOSION2POS
 564 => b"00000_0000_01_000000000000", -- load, gr0
 565 => b"00000_0000_00_000000000001", -- 1
 566 => b"00001_0000_10_010000101000", -- store, gr0, P2EXPLOSION2ACTIVE
 567 => b"00000_0000_01_000000000000", -- load, gr0
 568 => b"00000_0000_00_000000000010", -- 2
 569 => b"00001_0000_10_010000100111", -- store, gr0, P2EXPLOSION2TIME
 570 => b"00000_0000_00_010000110001", -- load, gr0, P2BOMBCOUNT
 571 => b"00011_0000_01_000000000000", -- sub, gr0
 572 => b"00000_0000_00_000000000001", -- 1
 573 => b"00001_0000_10_010000110001", -- store, gr0, P2BOMBCOUNT
 574 => b"00000_0100_00_010000100100", -- load, gr4, P2BOMB2POS
 575 => b"00100_0000_01_000000000000", -- jump
 576 => b"00000_0000_00_001001010011", -- EXPLODE
 577 => b"00000_0000_01_000000000000", -- load, gr0
 578 => b"00000_0000_00_000000000000", -- 0
 579 => b"00001_0000_10_010000101100", -- store, gr0, P2BOMB3ACTIVE
 580 => b"00000_0000_00_010000101010", -- load, gr0, P2BOMB3POS
 581 => b"00001_0000_10_010000101111", -- store, gr0, P2EXPLOSION3POS
 582 => b"00000_0000_01_000000000000", -- load, gr0
 583 => b"00000_0000_00_000000000001", -- 1
 584 => b"00001_0000_10_010000101110", -- store, gr0, P2EXPLOSION3ACTIVE
 585 => b"00000_0000_01_000000000000", -- load, gr0
 586 => b"00000_0000_00_000000000010", -- 2
 587 => b"00001_0000_10_010000101101", -- store, gr0, P2EXPLOSION3TIME
 588 => b"00000_0000_00_010000110001", -- load, gr0, P2BOMBCOUNT
 589 => b"00011_0000_01_000000000000", -- sub, gr0
 590 => b"00000_0000_00_000000000001", -- 1
 591 => b"00001_0000_10_010000110001", -- store, gr0, P2BOMBCOUNT
 592 => b"00000_0100_00_010000101010", -- load, gr4, P2BOMB3POS
 593 => b"00100_0000_01_000000000000", -- jump
 594 => b"00000_0000_00_001001010011", -- EXPLODE
 595 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 596 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 597 => b"00000_0011_00_010000111101", -- load, gr3, EXPLOSION
 598 => b"10000_0010_00_000000000000", -- tpoint, gr2
 599 => b"01110_0011_00_000000000000", -- twrite, gr3
 600 => b"00010_0010_01_000000000000", -- add, gr2
 601 => b"00000_0000_00_000000000001", -- 1
 602 => b"10000_0010_00_000000000000", -- tpoint, gr2
 603 => b"01111_0000_00_000000000000", -- tread, gr0
 604 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 605 => b"00110_0000_01_000000000000", -- beq
 606 => b"00000_0000_00_001001101000", -- EXPLODELEFT
 607 => b"01110_0011_00_000000000000", -- twrite, gr3
 608 => b"00010_0010_01_000000000000", -- add, gr2
 609 => b"00000_0000_00_000000000001", -- 1
 610 => b"10000_0010_00_000000000000", -- tpoint, gr2
 611 => b"01111_0000_00_000000000000", -- tread, gr0
 612 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 613 => b"00110_0000_01_000000000000", -- beq
 614 => b"00000_0000_00_001001101000", -- EXPLODELEFT
 615 => b"01110_0011_00_000000000000", -- twrite, gr3
 616 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 617 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 618 => b"00011_0010_01_000000000000", -- sub, gr2
 619 => b"00000_0000_00_000000000001", -- 1
 620 => b"10000_0010_00_000000000000", -- tpoint, gr2
 621 => b"01111_0000_00_000000000000", -- tread, gr0
 622 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 623 => b"00110_0000_01_000000000000", -- beq
 624 => b"00000_0000_00_001001111010", -- EXPLODEDOWN
 625 => b"01110_0011_00_000000000000", -- twrite, gr3
 626 => b"00011_0010_01_000000000000", -- sub, gr2
 627 => b"00000_0000_00_000000000001", -- 1
 628 => b"10000_0010_00_000000000000", -- tpoint, gr2
 629 => b"01111_0000_00_000000000000", -- tread, gr0
 630 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 631 => b"00110_0000_01_000000000000", -- beq
 632 => b"00000_0000_00_001001111010", -- EXPLODEDOWN
 633 => b"01110_0011_00_000000000000", -- twrite, gr3
 634 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 635 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 636 => b"00010_0010_01_000000000000", -- add, gr2
 637 => b"00000_0000_00_000000001111", -- 15
 638 => b"10000_0010_00_000000000000", -- tpoint, gr2
 639 => b"01111_0000_00_000000000000", -- tread, gr0
 640 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 641 => b"00110_0000_01_000000000000", -- beq
 642 => b"00000_0000_00_001010001100", -- EXPLODEUP
 643 => b"01110_0011_00_000000000000", -- twrite, gr3
 644 => b"00010_0010_01_000000000000", -- add, gr2
 645 => b"00000_0000_00_000000001111", -- 15
 646 => b"10000_0010_00_000000000000", -- tpoint, gr2
 647 => b"01111_0000_00_000000000000", -- tread, gr0
 648 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 649 => b"00110_0000_01_000000000000", -- beq
 650 => b"00000_0000_00_001010001100", -- EXPLODEUP
 651 => b"01110_0011_00_000000000000", -- twrite, gr3
 652 => b"00001_0100_10_010000110111", -- store, gr4, MOVE
 653 => b"00000_0010_00_010000110111", -- load, gr2, MOVE
 654 => b"00011_0010_01_000000000000", -- sub, gr2
 655 => b"00000_0000_00_000000001111", -- 15
 656 => b"10000_0010_00_000000000000", -- tpoint, gr2
 657 => b"01111_0000_00_000000000000", -- tread, gr0
 658 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 659 => b"00110_0000_01_000000000000", -- beq
 660 => b"00000_0000_00_000110010001", -- TICKBOMBS
 661 => b"01110_0011_00_000000000000", -- twrite, gr3
 662 => b"00011_0010_01_000000000000", -- sub, gr2
 663 => b"00000_0000_00_000000001111", -- 15
 664 => b"10000_0010_00_000000000000", -- tpoint, gr2
 665 => b"01111_0000_00_000000000000", -- tread, gr0
 666 => b"00011_0000_00_010000111011", -- sub, gr0, WALL
 667 => b"00110_0000_01_000000000000", -- beq
 668 => b"00000_0000_00_000110010001", -- TICKBOMBS
 669 => b"01110_0011_00_000000000000", -- twrite, gr3
 670 => b"00100_0000_01_000000000000", -- jump
 671 => b"00000_0000_00_000110010001", -- TICKBOMBS
 672 => b"10101_0000_01_000000000000", -- btn1
 673 => b"00000_0000_00_001010100110", -- BTN1
 674 => b"11010_0000_01_000000000000", -- btn2
 675 => b"00000_0000_00_001100000111", -- BTN2
 676 => b"00100_0000_01_000000000000", -- jump
 677 => b"00000_0000_00_000001101000", -- BUTTON_R
 678 => b"00000_0000_00_010000001010", -- load, gr0, P1DEAD
 679 => b"00011_0000_01_000000000000", -- sub, gr0
 680 => b"00000_0000_00_000000000001", -- 1
 681 => b"00110_0000_01_000000000000", -- beq
 682 => b"00000_0000_00_000000000000", -- INIT
 683 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMBCOUNT
 684 => b"00011_0000_00_010000110010", -- sub, gr0, MAXBOMBS
 685 => b"00110_0000_01_000000000000", -- beq
 686 => b"00000_0000_00_001010100010", -- BTN1_R
 687 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 688 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 689 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 690 => b"01000_0000_01_000000000000", -- mul, gr0
 691 => b"00000_0000_00_000000001111", -- 15
 692 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 693 => b"10000_0000_00_000000000000", -- tpoint, gr0
 694 => b"01111_0001_00_000000000000", -- tread, gr1
 695 => b"00011_0001_00_010000111110", -- sub, gr1, EGG
 696 => b"00110_0000_01_000000000000", -- beq
 697 => b"00000_0000_00_001010100010", -- BTN1_R
 698 => b"00000_0000_00_010000001110", -- load, gr0, P1BOMB1ACTIVE
 699 => b"00011_0000_01_000000000000", -- sub, gr0
 700 => b"00000_0000_00_000000000000", -- 0
 701 => b"00110_0000_01_000000000000", -- beq
 702 => b"00000_0000_00_001011010001", -- P1PLACEBOMB1
 703 => b"00000_0000_00_010000010100", -- load, gr0, P1BOMB2ACTIVE
 704 => b"00011_0000_01_000000000000", -- sub, gr0
 705 => b"00000_0000_00_000000000000", -- 0
 706 => b"00110_0000_01_000000000000", -- beq
 707 => b"00000_0000_00_001011100011", -- P1PLACEBOMB2
 708 => b"00000_0000_00_010000011010", -- load, gr0, P1BOMB3ACTIVE
 709 => b"00011_0000_01_000000000000", -- sub, gr0
 710 => b"00000_0000_00_000000000000", -- 0
 711 => b"00110_0000_01_000000000000", -- beq
 712 => b"00000_0000_00_001011110101", -- P1PLACEBOMB3
 713 => b"00100_0000_01_000000000000", -- jump
 714 => b"00000_0000_00_001010100010", -- BTN1_R
 715 => b"00000_0000_00_010000110000", -- load, gr0, P1BOMBCOUNT
 716 => b"00010_0000_01_000000000000", -- add, gr0
 717 => b"00000_0000_00_000000000001", -- 1
 718 => b"00001_0000_10_010000110000", -- store, gr0, P1BOMBCOUNT
 719 => b"00100_0000_01_000000000000", -- jump
 720 => b"00000_0000_00_001010100010", -- BTN1_R
 721 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 722 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 723 => b"00000_0011_00_010000110100", -- load, gr3, YPOS1
 724 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 725 => b"01000_0011_01_000000000000", -- mul, gr3
 726 => b"00000_0000_00_000000001111", -- 15
 727 => b"00010_0011_00_010000110011", -- add, gr3, XPOS1
 728 => b"10000_0011_00_000000000000", -- tpoint, gr3
 729 => b"01110_0010_00_000000000000", -- twrite, gr2
 730 => b"00000_0000_01_000000000000", -- load, gr0
 731 => b"00000_0000_00_000000000001", -- 1
 732 => b"00001_0000_10_010000001110", -- store, gr0, P1BOMB1ACTIVE
 733 => b"00001_0011_10_010000001100", -- store, gr3, P1BOMB1POS
 734 => b"00000_0000_01_000000000000", -- load, gr0
 735 => b"00000_0000_00_000000010000", -- 16
 736 => b"00001_0000_10_010000001101", -- store, gr0, P1BOMB1TIME
 737 => b"00100_0000_01_000000000000", -- jump
 738 => b"00000_0000_00_001011001011", -- P1INCREASEBOMBCOUNTER
 739 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 740 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 741 => b"00000_0011_00_010000110100", -- load, gr3, YPOS1
 742 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 743 => b"01000_0011_01_000000000000", -- mul, gr3
 744 => b"00000_0000_00_000000001111", -- 15
 745 => b"00010_0011_00_010000110011", -- add, gr3, XPOS1
 746 => b"10000_0011_00_000000000000", -- tpoint, gr3
 747 => b"01110_0010_00_000000000000", -- twrite, gr2
 748 => b"00000_0000_01_000000000000", -- load, gr0
 749 => b"00000_0000_00_000000000001", -- 1
 750 => b"00001_0000_10_010000010100", -- store, gr0, P1BOMB2ACTIVE
 751 => b"00001_0011_10_010000010010", -- store, gr3, P1BOMB2POS
 752 => b"00000_0000_01_000000000000", -- load, gr0
 753 => b"00000_0000_00_000000010000", -- 16
 754 => b"00001_0000_10_010000010011", -- store, gr0, P1BOMB2TIME
 755 => b"00100_0000_01_000000000000", -- jump
 756 => b"00000_0000_00_001011001011", -- P1INCREASEBOMBCOUNTER
 757 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 758 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 759 => b"00000_0011_00_010000110100", -- load, gr3, YPOS1
 760 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 761 => b"01000_0011_01_000000000000", -- mul, gr3
 762 => b"00000_0000_00_000000001111", -- 15
 763 => b"00010_0011_00_010000110011", -- add, gr3, XPOS1
 764 => b"10000_0011_00_000000000000", -- tpoint, gr3
 765 => b"01110_0010_00_000000000000", -- twrite, gr2
 766 => b"00000_0000_01_000000000000", -- load, gr0
 767 => b"00000_0000_00_000000000001", -- 1
 768 => b"00001_0000_10_010000011010", -- store, gr0, P1BOMB3ACTIVE
 769 => b"00001_0011_10_010000011000", -- store, gr3, P1BOMB3POS
 770 => b"00000_0000_01_000000000000", -- load, gr0
 771 => b"00000_0000_00_000000010000", -- 16
 772 => b"00001_0000_10_010000011001", -- store, gr0, P1BOMB3TIME
 773 => b"00100_0000_01_000000000000", -- jump
 774 => b"00000_0000_00_001011001011", -- P1INCREASEBOMBCOUNTER
 775 => b"00000_0000_00_010000001011", -- load, gr0, P2DEAD
 776 => b"00011_0000_01_000000000000", -- sub, gr0
 777 => b"00000_0000_00_000000000001", -- 1
 778 => b"00110_0000_01_000000000000", -- beq
 779 => b"00000_0000_00_000000000000", -- INIT
 780 => b"00000_0000_00_010000110001", -- load, gr0, P2BOMBCOUNT
 781 => b"00011_0000_00_010000110010", -- sub, gr0, MAXBOMBS
 782 => b"00110_0000_01_000000000000", -- beq
 783 => b"00000_0000_00_001010100100", -- BTN2_R
 784 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 785 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 786 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
 787 => b"01000_0000_01_000000000000", -- mul, gr0
 788 => b"00000_0000_00_000000001111", -- 15
 789 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
 790 => b"10000_0000_00_000000000000", -- tpoint, gr0
 791 => b"01111_0001_00_000000000000", -- tread, gr1
 792 => b"00011_0001_00_010000111110", -- sub, gr1, EGG
 793 => b"00110_0000_01_000000000000", -- beq
 794 => b"00000_0000_00_001010100100", -- BTN2_R
 795 => b"00000_0000_00_010000100000", -- load, gr0, P2BOMB1ACTIVE
 796 => b"00011_0000_01_000000000000", -- sub, gr0
 797 => b"00000_0000_00_000000000000", -- 0
 798 => b"00110_0000_01_000000000000", -- beq
 799 => b"00000_0000_00_001100110000", -- P2PLACEBOMB1
 800 => b"00000_0000_00_010000100110", -- load, gr0, P2BOMB2ACTIVE
 801 => b"00011_0000_01_000000000000", -- sub, gr0
 802 => b"00000_0000_00_000000000000", -- 0
 803 => b"00110_0000_01_000000000000", -- beq
 804 => b"00000_0000_00_001101000010", -- P2PLACEBOMB2
 805 => b"00000_0000_00_010000101100", -- load, gr0, P2BOMB3ACTIVE
 806 => b"00011_0000_01_000000000000", -- sub, gr0
 807 => b"00000_0000_00_000000000000", -- 0
 808 => b"00110_0000_01_000000000000", -- beq
 809 => b"00000_0000_00_001101010100", -- P2PLACEBOMB3
 810 => b"00000_0000_00_010000110001", -- load, gr0, P2BOMBCOUNT
 811 => b"00010_0000_01_000000000000", -- add, gr0
 812 => b"00000_0000_00_000000000001", -- 1
 813 => b"00001_0000_10_010000110001", -- store, gr0, P2BOMBCOUNT
 814 => b"00100_0000_01_000000000000", -- jump
 815 => b"00000_0000_00_001010100100", -- BTN2_R
 816 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 817 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 818 => b"00000_0011_00_010000110110", -- load, gr3, YPOS2
 819 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 820 => b"01000_0011_01_000000000000", -- mul, gr3
 821 => b"00000_0000_00_000000001111", -- 15
 822 => b"00010_0011_00_010000110101", -- add, gr3, XPOS2
 823 => b"10000_0011_00_000000000000", -- tpoint, gr3
 824 => b"01110_0010_00_000000000000", -- twrite, gr2
 825 => b"00000_0000_01_000000000000", -- load, gr0
 826 => b"00000_0000_00_000000000001", -- 1
 827 => b"00001_0000_10_010000100000", -- store, gr0, P2BOMB1ACTIVE
 828 => b"00001_0011_10_010000011110", -- store, gr3, P2BOMB1POS
 829 => b"00000_0000_01_000000000000", -- load, gr0
 830 => b"00000_0000_00_000000010000", -- 16
 831 => b"00001_0000_10_010000011111", -- store, gr0, P2BOMB1TIME
 832 => b"00100_0000_01_000000000000", -- jump
 833 => b"00000_0000_00_001100101010", -- P2INCREASEBOMBCOUNTER
 834 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 835 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 836 => b"00000_0011_00_010000110110", -- load, gr3, YPOS2
 837 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 838 => b"01000_0011_01_000000000000", -- mul, gr3
 839 => b"00000_0000_00_000000001111", -- 15
 840 => b"00010_0011_00_010000110101", -- add, gr3, XPOS2
 841 => b"10000_0011_00_000000000000", -- tpoint, gr3
 842 => b"01110_0010_00_000000000000", -- twrite, gr2
 843 => b"00000_0000_01_000000000000", -- load, gr0
 844 => b"00000_0000_00_000000000001", -- 1
 845 => b"00001_0000_10_010000100110", -- store, gr0, P2BOMB2ACTIVE
 846 => b"00001_0011_10_010000100100", -- store, gr3, P2BOMB2POS
 847 => b"00000_0000_01_000000000000", -- load, gr0
 848 => b"00000_0000_00_000000010000", -- 16
 849 => b"00001_0000_10_010000100101", -- store, gr0, P2BOMB2TIME
 850 => b"00100_0000_01_000000000000", -- jump
 851 => b"00000_0000_00_001100101010", -- P2INCREASEBOMBCOUNTER
 852 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 853 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 854 => b"00000_0011_00_010000110110", -- load, gr3, YPOS2
 855 => b"00000_0010_00_010000111110", -- load, gr2, EGG
 856 => b"01000_0011_01_000000000000", -- mul, gr3
 857 => b"00000_0000_00_000000001111", -- 15
 858 => b"00010_0011_00_010000110101", -- add, gr3, XPOS2
 859 => b"10000_0011_00_000000000000", -- tpoint, gr3
 860 => b"01110_0010_00_000000000000", -- twrite, gr2
 861 => b"00000_0000_01_000000000000", -- load, gr0
 862 => b"00000_0000_00_000000000001", -- 1
 863 => b"00001_0000_10_010000101100", -- store, gr0, P2BOMB3ACTIVE
 864 => b"00001_0011_10_010000101010", -- store, gr3, P2BOMB3POS
 865 => b"00000_0000_01_000000000000", -- load, gr0
 866 => b"00000_0000_00_000000010000", -- 16
 867 => b"00001_0000_10_010000101011", -- store, gr0, P2BOMB3TIME
 868 => b"00100_0000_01_000000000000", -- jump
 869 => b"00000_0000_00_001100101010", -- P2INCREASEBOMBCOUNTER
 870 => b"00000_0000_00_010000001010", -- load, gr0, P1DEAD
 871 => b"00011_0000_01_000000000000", -- sub, gr0
 872 => b"00000_0000_00_000000000001", -- 1
 873 => b"00110_0000_01_000000000000", -- beq
 874 => b"00000_0000_00_001101110011", -- J2
 875 => b"10001_0000_01_000000000000", -- joy1r
 876 => b"00000_0000_00_001110000010", -- P1R
 877 => b"10011_0000_01_000000000000", -- joy1l
 878 => b"00000_0000_00_001110100100", -- P1L
 879 => b"10010_0000_01_000000000000", -- joy1u
 880 => b"00000_0000_00_001110010011", -- P1U
 881 => b"10100_0000_01_000000000000", -- joy1d
 882 => b"00000_0000_00_001110110101", -- P1D
 883 => b"00000_0000_00_010000001011", -- load, gr0, P2DEAD
 884 => b"00011_0000_01_000000000000", -- sub, gr0
 885 => b"00000_0000_00_000000000001", -- 1
 886 => b"00110_0000_01_000000000000", -- beq
 887 => b"00000_0000_00_000001100110", -- CONTROL_R
 888 => b"10110_0000_01_000000000000", -- joy2r
 889 => b"00000_0000_00_001111000110", -- P2R
 890 => b"11000_0000_01_000000000000", -- joy2l
 891 => b"00000_0000_00_001111101000", -- P2L
 892 => b"10111_0000_01_000000000000", -- joy2u
 893 => b"00000_0000_00_001111010111", -- P2U
 894 => b"11001_0000_01_000000000000", -- joy2d
 895 => b"00000_0000_00_001111111001", -- P2D
 896 => b"00100_0000_01_000000000000", -- jump
 897 => b"00000_0000_00_000001100110", -- CONTROL_R
 898 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 899 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 900 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 901 => b"01000_0000_01_000000000000", -- mul, gr0
 902 => b"00000_0000_00_000000001111", -- 15
 903 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 904 => b"00010_0000_01_000000000000", -- add, gr0
 905 => b"00000_0000_00_000000000001", -- 1
 906 => b"10000_0000_00_000000000000", -- tpoint, gr0
 907 => b"01111_0001_00_000000000000", -- tread, gr1
 908 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 909 => b"00111_0000_01_000000000000", -- bne
 910 => b"00000_0000_00_001101101111", -- J1
 911 => b"00010_1100_01_000000000000", -- add, gr12
 912 => b"00000_0000_00_000000000001", -- 1
 913 => b"00100_0000_01_000000000000", -- jump
 914 => b"00000_0000_00_001101101111", -- J1
 915 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 916 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 917 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 918 => b"00011_0000_01_000000000000", -- sub, gr0
 919 => b"00000_0000_00_000000000001", -- 1
 920 => b"01000_0000_01_000000000000", -- mul, gr0
 921 => b"00000_0000_00_000000001111", -- 15
 922 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 923 => b"10000_0000_00_000000000000", -- tpoint, gr0
 924 => b"01111_0001_00_000000000000", -- tread, gr1
 925 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 926 => b"00111_0000_01_000000000000", -- bne
 927 => b"00000_0000_00_001101110011", -- J2
 928 => b"00011_1101_01_000000000000", -- sub, gr13
 929 => b"00000_0000_00_000000000001", -- 1
 930 => b"00100_0000_01_000000000000", -- jump
 931 => b"00000_0000_00_001101110011", -- J2
 932 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 933 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 934 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 935 => b"01000_0000_01_000000000000", -- mul, gr0
 936 => b"00000_0000_00_000000001111", -- 15
 937 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 938 => b"00011_0000_01_000000000000", -- sub, gr0
 939 => b"00000_0000_00_000000000001", -- 1
 940 => b"10000_0000_00_000000000000", -- tpoint, gr0
 941 => b"01111_0001_00_000000000000", -- tread, gr1
 942 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 943 => b"00111_0000_01_000000000000", -- bne
 944 => b"00000_0000_00_001101101111", -- J1
 945 => b"00011_1100_01_000000000000", -- sub, gr12
 946 => b"00000_0000_00_000000000001", -- 1
 947 => b"00100_0000_01_000000000000", -- jump
 948 => b"00000_0000_00_001101101111", -- J1
 949 => b"00001_1100_10_010000110011", -- store, gr12, XPOS1
 950 => b"00001_1101_10_010000110100", -- store, gr13, YPOS1
 951 => b"00000_0000_00_010000110100", -- load, gr0, YPOS1
 952 => b"00010_0000_01_000000000000", -- add, gr0
 953 => b"00000_0000_00_000000000001", -- 1
 954 => b"01000_0000_01_000000000000", -- mul, gr0
 955 => b"00000_0000_00_000000001111", -- 15
 956 => b"00010_0000_00_010000110011", -- add, gr0, XPOS1
 957 => b"10000_0000_00_000000000000", -- tpoint, gr0
 958 => b"01111_0001_00_000000000000", -- tread, gr1
 959 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 960 => b"00111_0000_01_000000000000", -- bne
 961 => b"00000_0000_00_001101110011", -- J2
 962 => b"00010_1101_01_000000000000", -- add, gr13
 963 => b"00000_0000_00_000000000001", -- 1
 964 => b"00100_0000_01_000000000000", -- jump
 965 => b"00000_0000_00_001101110011", -- J2
 966 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 967 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 968 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
 969 => b"01000_0000_01_000000000000", -- mul, gr0
 970 => b"00000_0000_00_000000001111", -- 15
 971 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
 972 => b"00010_0000_01_000000000000", -- add, gr0
 973 => b"00000_0000_00_000000000001", -- 1
 974 => b"10000_0000_00_000000000000", -- tpoint, gr0
 975 => b"01111_0001_00_000000000000", -- tread, gr1
 976 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 977 => b"00111_0000_01_000000000000", -- bne
 978 => b"00000_0000_00_001101111100", -- J3
 979 => b"00010_1110_01_000000000000", -- add, gr14
 980 => b"00000_0000_00_000000000001", -- 1
 981 => b"00100_0000_01_000000000000", -- jump
 982 => b"00000_0000_00_001101111100", -- J3
 983 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
 984 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
 985 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
 986 => b"00011_0000_01_000000000000", -- sub, gr0
 987 => b"00000_0000_00_000000000001", -- 1
 988 => b"01000_0000_01_000000000000", -- mul, gr0
 989 => b"00000_0000_00_000000001111", -- 15
 990 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
 991 => b"10000_0000_00_000000000000", -- tpoint, gr0
 992 => b"01111_0001_00_000000000000", -- tread, gr1
 993 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
 994 => b"00111_0000_01_000000000000", -- bne
 995 => b"00000_0000_00_000001100110", -- CONTROL_R
 996 => b"00011_1111_01_000000000000", -- sub, gr15
 997 => b"00000_0000_00_000000000001", -- 1
 998 => b"00100_0000_01_000000000000", -- jump
 999 => b"00000_0000_00_000001100110", -- CONTROL_R
1000 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
1001 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
1002 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
1003 => b"01000_0000_01_000000000000", -- mul, gr0
1004 => b"00000_0000_00_000000001111", -- 15
1005 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
1006 => b"00011_0000_01_000000000000", -- sub, gr0
1007 => b"00000_0000_00_000000000001", -- 1
1008 => b"10000_0000_00_000000000000", -- tpoint, gr0
1009 => b"01111_0001_00_000000000000", -- tread, gr1
1010 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
1011 => b"00111_0000_01_000000000000", -- bne
1012 => b"00000_0000_00_001101111100", -- J3
1013 => b"00011_1110_01_000000000000", -- sub, gr14
1014 => b"00000_0000_00_000000000001", -- 1
1015 => b"00100_0000_01_000000000000", -- jump
1016 => b"00000_0000_00_001101111100", -- J3
1017 => b"00001_1110_10_010000110101", -- store, gr14, XPOS2
1018 => b"00001_1111_10_010000110110", -- store, gr15, YPOS2
1019 => b"00000_0000_00_010000110110", -- load, gr0, YPOS2
1020 => b"00010_0000_01_000000000000", -- add, gr0
1021 => b"00000_0000_00_000000000001", -- 1
1022 => b"01000_0000_01_000000000000", -- mul, gr0
1023 => b"00000_0000_00_000000001111", -- 15
1024 => b"00010_0000_00_010000110101", -- add, gr0, XPOS2
1025 => b"10000_0000_00_000000000000", -- tpoint, gr0
1026 => b"01111_0001_00_000000000000", -- tread, gr1
1027 => b"00011_0001_00_010000111010", -- sub, gr1, GRASS
1028 => b"00111_0000_01_000000000000", -- bne
1029 => b"00000_0000_00_000001100110", -- CONTROL_R
1030 => b"00010_1111_01_000000000000", -- add, gr15
1031 => b"00000_0000_00_000000000001", -- 1
1032 => b"00100_0000_01_000000000000", -- jump
1033 => b"00000_0000_00_000001100110", -- CONTROL_R
1034 => b"00000_0000_00_000000000000", -- 0
1035 => b"00000_0000_00_000000000000", -- 0
1036 => b"00000_0000_00_000000000000", -- 0
1037 => b"00000_0000_00_000000000000", -- 0
1038 => b"00000_0000_00_000000000000", -- 0
1039 => b"00000_0000_00_000000000000", -- 0
1040 => b"00000_0000_00_000000000000", -- 0
1041 => b"00000_0000_00_000000000000", -- 0
1042 => b"00000_0000_00_000000000000", -- 0
1043 => b"00000_0000_00_000000000000", -- 0
1044 => b"00000_0000_00_000000000000", -- 0
1045 => b"00000_0000_00_000000000000", -- 0
1046 => b"00000_0000_00_000000000000", -- 0
1047 => b"00000_0000_00_000000000000", -- 0
1048 => b"00000_0000_00_000000000000", -- 0
1049 => b"00000_0000_00_000000000000", -- 0
1050 => b"00000_0000_00_000000000000", -- 0
1051 => b"00000_0000_00_000000000000", -- 0
1052 => b"00000_0000_00_000000000000", -- 0
1053 => b"00000_0000_00_000000000000", -- 0
1054 => b"00000_0000_00_000000000000", -- 0
1055 => b"00000_0000_00_000000000000", -- 0
1056 => b"00000_0000_00_000000000000", -- 0
1057 => b"00000_0000_00_000000000000", -- 0
1058 => b"00000_0000_00_000000000000", -- 0
1059 => b"00000_0000_00_000000000000", -- 0
1060 => b"00000_0000_00_000000000000", -- 0
1061 => b"00000_0000_00_000000000000", -- 0
1062 => b"00000_0000_00_000000000000", -- 0
1063 => b"00000_0000_00_000000000000", -- 0
1064 => b"00000_0000_00_000000000000", -- 0
1065 => b"00000_0000_00_000000000000", -- 0
1066 => b"00000_0000_00_000000000000", -- 0
1067 => b"00000_0000_00_000000000000", -- 0
1068 => b"00000_0000_00_000000000000", -- 0
1069 => b"00000_0000_00_000000000000", -- 0
1070 => b"00000_0000_00_000000000000", -- 0
1071 => b"00000_0000_00_000000000000", -- 0
1072 => b"00000_0000_00_000000000000", -- 0
1073 => b"00000_0000_00_000000000000", -- 0
1074 => b"00000_0000_00_000000000011", -- 3
1075 => b"00000_0000_00_000000000000", -- 0
1076 => b"00000_0000_00_000000000000", -- 0
1077 => b"00000_0000_00_000000000000", -- 0
1078 => b"00000_0000_00_000000000000", -- 0
1079 => b"00000_0000_00_000000000000", -- 0
1080 => b"00000_0000_00_000000000000", -- 0
1081 => b"00000_0000_00_000000000000", -- 0
1082 => b"00000_0000_00_000000000000", -- 0
1083 => b"00000_0000_00_000000000001", -- 1
1084 => b"00000_0000_00_000000000010", -- 2
1085 => b"00000_0000_00_000000000011", -- 3
1086 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
