library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_001010011100", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000111100000", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011010001", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00000_0000_00_001100111110", -- load, gr0, P1EXPLOSION1ACTIVE
  11 => b"00011_0000_01_000000000000", -- sub, gr0
  12 => b"00000_0000_00_000000000001", -- 1
  13 => b"00111_0000_01_000000000000", -- bne
  14 => b"00000_0000_00_000000011000", -- P1EXPLOSION2
  15 => b"00000_0000_00_001100111101", -- load, gr0, P1EXPLOSION1TIME
  16 => b"00011_0000_01_000000000000", -- sub, gr0
  17 => b"00000_0000_00_000000000001", -- 1
  18 => b"00001_0000_10_001100111101", -- store, gr0, P1EXPLOSION1TIME
  19 => b"00000_0000_01_000000000000", -- load, gr0
  20 => b"00000_0000_00_000000000000", -- 0
  21 => b"00011_0000_00_001100111101", -- sub, gr0, P1EXPLOSION1TIME
  22 => b"00110_0000_01_000000000000", -- beq
  23 => b"00000_0000_00_000001100000", -- P1EXPLOSION1FADE
  24 => b"00000_0000_00_001101000100", -- load, gr0, P1EXPLOSION2ACTIVE
  25 => b"00011_0000_01_000000000000", -- sub, gr0
  26 => b"00000_0000_00_000000000001", -- 1
  27 => b"00111_0000_01_000000000000", -- bne
  28 => b"00000_0000_00_000000100110", -- P1EXPLOSION3
  29 => b"00000_0000_00_001101000011", -- load, gr0, P1EXPLOSION2TIME
  30 => b"00011_0000_01_000000000000", -- sub, gr0
  31 => b"00000_0000_00_000000000001", -- 1
  32 => b"00001_0000_10_001101000011", -- store, gr0, P1EXPLOSION2TIME
  33 => b"00000_0000_01_000000000000", -- load, gr0
  34 => b"00000_0000_00_000000000000", -- 0
  35 => b"00011_0000_00_001101000011", -- sub, gr0, P1EXPLOSION2TIME
  36 => b"00110_0000_01_000000000000", -- beq
  37 => b"00000_0000_00_000001100110", -- P1EXPLOSION2FADE
  38 => b"00000_0000_00_001101001010", -- load, gr0, P1EXPLOSION3ACTIVE
  39 => b"00011_0000_01_000000000000", -- sub, gr0
  40 => b"00000_0000_00_000000000001", -- 1
  41 => b"00111_0000_01_000000000000", -- bne
  42 => b"00000_0000_00_000000110100", -- P2EXPLOSION1
  43 => b"00000_0000_00_001101001001", -- load, gr0, P1EXPLOSION3TIME
  44 => b"00011_0000_01_000000000000", -- sub, gr0
  45 => b"00000_0000_00_000000000001", -- 1
  46 => b"00001_0000_10_001101001001", -- store, gr0, P1EXPLOSION3TIME
  47 => b"00000_0000_01_000000000000", -- load, gr0
  48 => b"00000_0000_00_000000000000", -- 0
  49 => b"00011_0000_00_001101001001", -- sub, gr0, P1EXPLOSION3TIME
  50 => b"00110_0000_01_000000000000", -- beq
  51 => b"00000_0000_00_000001101100", -- P1EXPLOSION3FADE
  52 => b"00000_0000_00_001101010000", -- load, gr0, P2EXPLOSION1ACTIVE
  53 => b"00011_0000_01_000000000000", -- sub, gr0
  54 => b"00000_0000_00_000000000001", -- 1
  55 => b"00111_0000_01_000000000000", -- bne
  56 => b"00000_0000_00_000001000010", -- P2EXPLOSION2
  57 => b"00000_0000_00_001101001111", -- load, gr0, P2EXPLOSION1TIME
  58 => b"00011_0000_01_000000000000", -- sub, gr0
  59 => b"00000_0000_00_000000000001", -- 1
  60 => b"00001_0000_10_001101001111", -- store, gr0, P2EXPLOSION1TIME
  61 => b"00000_0000_01_000000000000", -- load, gr0
  62 => b"00000_0000_00_000000000000", -- 0
  63 => b"00011_0000_00_001101001111", -- sub, gr0, P2EXPLOSION1TIME
  64 => b"00110_0000_01_000000000000", -- beq
  65 => b"00000_0000_00_000001110010", -- P2EXPLOSION1FADE
  66 => b"00000_0000_00_001101010110", -- load, gr0, P2EXPLOSION2ACTIVE
  67 => b"00011_0000_01_000000000000", -- sub, gr0
  68 => b"00000_0000_00_000000000001", -- 1
  69 => b"00111_0000_01_000000000000", -- bne
  70 => b"00000_0000_00_000001010000", -- P2EXPLOSION3
  71 => b"00000_0000_00_001101010101", -- load, gr0, P2EXPLOSION2TIME
  72 => b"00011_0000_01_000000000000", -- sub, gr0
  73 => b"00000_0000_00_000000000001", -- 1
  74 => b"00001_0000_10_001101010101", -- store, gr0, P2EXPLOSION2TIME
  75 => b"00000_0000_01_000000000000", -- load, gr0
  76 => b"00000_0000_00_000000000000", -- 0
  77 => b"00011_0000_00_001101010101", -- sub, gr0, P2EXPLOSION2TIME
  78 => b"00110_0000_01_000000000000", -- beq
  79 => b"00000_0000_00_000001111000", -- P2EXPLOSION2FADE
  80 => b"00000_0000_00_001101011100", -- load, gr0, P2EXPLOSION3ACTIVE
  81 => b"00011_0000_01_000000000000", -- sub, gr0
  82 => b"00000_0000_00_000000000001", -- 1
  83 => b"00111_0000_01_000000000000", -- bne
  84 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  85 => b"00000_0000_00_001101011011", -- load, gr0, P2EXPLOSION3TIME
  86 => b"00011_0000_01_000000000000", -- sub, gr0
  87 => b"00000_0000_00_000000000001", -- 1
  88 => b"00001_0000_10_001101011011", -- store, gr0, P2EXPLOSION3TIME
  89 => b"00000_0000_01_000000000000", -- load, gr0
  90 => b"00000_0000_00_000000000000", -- 0
  91 => b"00011_0000_00_001101011011", -- sub, gr0, P2EXPLOSION3TIME
  92 => b"00110_0000_01_000000000000", -- beq
  93 => b"00000_0000_00_000001111110", -- P2EXPLOSION3FADE
  94 => b"00100_0000_01_000000000000", -- jump
  95 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  96 => b"00000_0000_01_000000000000", -- load, gr0
  97 => b"00000_0000_00_000000000000", -- 0
  98 => b"00001_0000_10_001100111110", -- store, gr0, P1EXPLOSION1ACTIVE
  99 => b"00000_0100_00_001100111111", -- load, gr4, P1EXPLOSION1POS
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 102 => b"00000_0000_01_000000000000", -- load, gr0
 103 => b"00000_0000_00_000000000000", -- 0
 104 => b"00001_0000_10_001101000100", -- store, gr0, P1EXPLOSION2ACTIVE
 105 => b"00000_0100_00_001101000101", -- load, gr4, P1EXPLOSION2POS
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 108 => b"00000_0000_01_000000000000", -- load, gr0
 109 => b"00000_0000_00_000000000000", -- 0
 110 => b"00001_0000_10_001101001010", -- store, gr0, P1EXPLOSION3ACTIVE
 111 => b"00000_0100_00_001101001011", -- load, gr4, P1EXPLOSION3POS
 112 => b"00100_0000_01_000000000000", -- jump
 113 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 114 => b"00000_0000_01_000000000000", -- load, gr0
 115 => b"00000_0000_00_000000000000", -- 0
 116 => b"00001_0000_10_001101010000", -- store, gr0, P2EXPLOSION1ACTIVE
 117 => b"00000_0100_00_001101010001", -- load, gr4, P2EXPLOSION1POS
 118 => b"00100_0000_01_000000000000", -- jump
 119 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001101010110", -- store, gr0, P2EXPLOSION2ACTIVE
 123 => b"00000_0100_00_001101010111", -- load, gr4, P2EXPLOSION2POS
 124 => b"00100_0000_01_000000000000", -- jump
 125 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 126 => b"00000_0000_01_000000000000", -- load, gr0
 127 => b"00000_0000_00_000000000000", -- 0
 128 => b"00001_0000_10_001101011100", -- store, gr0, P2EXPLOSION3ACTIVE
 129 => b"00000_0100_00_001101011101", -- load, gr4, P2EXPLOSION3POS
 130 => b"00100_0000_01_000000000000", -- jump
 131 => b"00000_0000_00_000010000100", -- FADEEXPLOSION
 132 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 133 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 134 => b"00000_0011_00_001101101000", -- load, gr3, GRASS
 135 => b"10000_0010_00_000000000000", -- tpoint, gr2
 136 => b"01110_0011_00_000000000000", -- twrite, gr3
 137 => b"00010_0010_01_000000000000", -- add, gr2
 138 => b"00000_0000_00_000000000001", -- 1
 139 => b"10000_0010_00_000000000000", -- tpoint, gr2
 140 => b"01111_0000_00_000000000000", -- tread, gr0
 141 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 142 => b"00111_0000_01_000000000000", -- bne
 143 => b"00000_0000_00_000010011001", -- FADELEFT
 144 => b"01110_0011_00_000000000000", -- twrite, gr3
 145 => b"00010_0010_01_000000000000", -- add, gr2
 146 => b"00000_0000_00_000000000001", -- 1
 147 => b"10000_0010_00_000000000000", -- tpoint, gr2
 148 => b"01111_0000_00_000000000000", -- tread, gr0
 149 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 150 => b"00111_0000_01_000000000000", -- bne
 151 => b"00000_0000_00_000010011001", -- FADELEFT
 152 => b"01110_0011_00_000000000000", -- twrite, gr3
 153 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 154 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 155 => b"00011_0010_01_000000000000", -- sub, gr2
 156 => b"00000_0000_00_000000000001", -- 1
 157 => b"10000_0010_00_000000000000", -- tpoint, gr2
 158 => b"01111_0000_00_000000000000", -- tread, gr0
 159 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 160 => b"00111_0000_01_000000000000", -- bne
 161 => b"00000_0000_00_000010101011", -- FADEDOWN
 162 => b"01110_0011_00_000000000000", -- twrite, gr3
 163 => b"00011_0010_01_000000000000", -- sub, gr2
 164 => b"00000_0000_00_000000000001", -- 1
 165 => b"10000_0010_00_000000000000", -- tpoint, gr2
 166 => b"01111_0000_00_000000000000", -- tread, gr0
 167 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 168 => b"00111_0000_01_000000000000", -- bne
 169 => b"00000_0000_00_000010101011", -- FADEDOWN
 170 => b"01110_0011_00_000000000000", -- twrite, gr3
 171 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 172 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 173 => b"00010_0010_01_000000000000", -- add, gr2
 174 => b"00000_0000_00_000000001111", -- 15
 175 => b"10000_0010_00_000000000000", -- tpoint, gr2
 176 => b"01111_0000_00_000000000000", -- tread, gr0
 177 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 178 => b"00111_0000_01_000000000000", -- bne
 179 => b"00000_0000_00_000010111101", -- FADEUP
 180 => b"01110_0011_00_000000000000", -- twrite, gr3
 181 => b"00010_0010_01_000000000000", -- add, gr2
 182 => b"00000_0000_00_000000001111", -- 15
 183 => b"10000_0010_00_000000000000", -- tpoint, gr2
 184 => b"01111_0000_00_000000000000", -- tread, gr0
 185 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 186 => b"00111_0000_01_000000000000", -- bne
 187 => b"00000_0000_00_000010111101", -- FADEUP
 188 => b"01110_0011_00_000000000000", -- twrite, gr3
 189 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 190 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 191 => b"00011_0010_01_000000000000", -- sub, gr2
 192 => b"00000_0000_00_000000001111", -- 15
 193 => b"10000_0010_00_000000000000", -- tpoint, gr2
 194 => b"01111_0000_00_000000000000", -- tread, gr0
 195 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 196 => b"00111_0000_01_000000000000", -- bne
 197 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
 198 => b"01110_0011_00_000000000000", -- twrite, gr3
 199 => b"00011_0010_01_000000000000", -- sub, gr2
 200 => b"00000_0000_00_000000001111", -- 15
 201 => b"10000_0010_00_000000000000", -- tpoint, gr2
 202 => b"01111_0000_00_000000000000", -- tread, gr0
 203 => b"00011_0000_00_001101101011", -- sub, gr0, EXPLOSION
 204 => b"00111_0000_01_000000000000", -- bne
 205 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
 206 => b"01110_0011_00_000000000000", -- twrite, gr3
 207 => b"00100_0000_01_000000000000", -- jump
 208 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
 209 => b"00000_0000_00_001100111100", -- load, gr0, P1BOMB1ACTIVE
 210 => b"00011_0000_01_000000000000", -- sub, gr0
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00111_0000_01_000000000000", -- bne
 213 => b"00000_0000_00_000011011111", -- P1BOMB2
 214 => b"00000_0000_00_001100111011", -- load, gr0, P1BOMB1TIME
 215 => b"00011_0000_01_000000000000", -- sub, gr0
 216 => b"00000_0000_00_000000000001", -- 1
 217 => b"00001_0000_10_001100111011", -- store, gr0, P1BOMB1TIME
 218 => b"00000_0000_01_000000000000", -- load, gr0
 219 => b"00000_0000_00_000000000000", -- 0
 220 => b"00011_0000_00_001100111011", -- sub, gr0, P1BOMB1TIME
 221 => b"00110_0000_01_000000000000", -- beq
 222 => b"00000_0000_00_000100100111", -- P1EXPLOSION1INIT
 223 => b"00000_0000_00_001101000010", -- load, gr0, P1BOMB2ACTIVE
 224 => b"00011_0000_01_000000000000", -- sub, gr0
 225 => b"00000_0000_00_000000000001", -- 1
 226 => b"00111_0000_01_000000000000", -- bne
 227 => b"00000_0000_00_000011101101", -- P1BOMB3
 228 => b"00000_0000_00_001101000001", -- load, gr0, P1BOMB2TIME
 229 => b"00011_0000_01_000000000000", -- sub, gr0
 230 => b"00000_0000_00_000000000001", -- 1
 231 => b"00001_0000_10_001101000001", -- store, gr0, P1BOMB2TIME
 232 => b"00000_0000_01_000000000000", -- load, gr0
 233 => b"00000_0000_00_000000000000", -- 0
 234 => b"00011_0000_00_001101000001", -- sub, gr0, P1BOMB2TIME
 235 => b"00110_0000_01_000000000000", -- beq
 236 => b"00000_0000_00_000100111001", -- P1EXPLOSION2INIT
 237 => b"00000_0000_00_001101001000", -- load, gr0, P1BOMB3ACTIVE
 238 => b"00011_0000_01_000000000000", -- sub, gr0
 239 => b"00000_0000_00_000000000001", -- 1
 240 => b"00111_0000_01_000000000000", -- bne
 241 => b"00000_0000_00_000011111011", -- P2BOMB1
 242 => b"00000_0000_00_001101000111", -- load, gr0, P1BOMB3TIME
 243 => b"00011_0000_01_000000000000", -- sub, gr0
 244 => b"00000_0000_00_000000000001", -- 1
 245 => b"00001_0000_10_001101000111", -- store, gr0, P1BOMB3TIME
 246 => b"00000_0000_01_000000000000", -- load, gr0
 247 => b"00000_0000_00_000000000000", -- 0
 248 => b"00011_0000_00_001101000111", -- sub, gr0, P1BOMB3TIME
 249 => b"00110_0000_01_000000000000", -- beq
 250 => b"00000_0000_00_000101001011", -- P1EXPLOSION3INIT
 251 => b"00000_0000_00_001101001110", -- load, gr0, P2BOMB1ACTIVE
 252 => b"00011_0000_01_000000000000", -- sub, gr0
 253 => b"00000_0000_00_000000000001", -- 1
 254 => b"00111_0000_01_000000000000", -- bne
 255 => b"00000_0000_00_000100001001", -- P2BOMB2
 256 => b"00000_0000_00_001101001101", -- load, gr0, P2BOMB1TIME
 257 => b"00011_0000_01_000000000000", -- sub, gr0
 258 => b"00000_0000_00_000000000001", -- 1
 259 => b"00001_0000_10_001101001101", -- store, gr0, P2BOMB1TIME
 260 => b"00000_0000_01_000000000000", -- load, gr0
 261 => b"00000_0000_00_000000000000", -- 0
 262 => b"00011_0000_00_001101001101", -- sub, gr0, P2BOMB1TIME
 263 => b"00110_0000_01_000000000000", -- beq
 264 => b"00000_0000_00_000101011101", -- P2EXPLOSION1INIT
 265 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMB2ACTIVE
 266 => b"00011_0000_01_000000000000", -- sub, gr0
 267 => b"00000_0000_00_000000000001", -- 1
 268 => b"00111_0000_01_000000000000", -- bne
 269 => b"00000_0000_00_000100010111", -- P2BOMB3
 270 => b"00000_0000_00_001101010011", -- load, gr0, P2BOMB2TIME
 271 => b"00011_0000_01_000000000000", -- sub, gr0
 272 => b"00000_0000_00_000000000001", -- 1
 273 => b"00001_0000_10_001101010011", -- store, gr0, P2BOMB2TIME
 274 => b"00000_0000_01_000000000000", -- load, gr0
 275 => b"00000_0000_00_000000000000", -- 0
 276 => b"00011_0000_00_001101010011", -- sub, gr0, P2BOMB2TIME
 277 => b"00110_0000_01_000000000000", -- beq
 278 => b"00000_0000_00_000101101111", -- P2EXPLOSION2INIT
 279 => b"00000_0000_00_001101011010", -- load, gr0, P2BOMB3ACTIVE
 280 => b"00011_0000_01_000000000000", -- sub, gr0
 281 => b"00000_0000_00_000000000001", -- 1
 282 => b"00111_0000_01_000000000000", -- bne
 283 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 284 => b"00000_0000_00_001101011001", -- load, gr0, P2BOMB3TIME
 285 => b"00011_0000_01_000000000000", -- sub, gr0
 286 => b"00000_0000_00_000000000001", -- 1
 287 => b"00001_0000_10_001101011001", -- store, gr0, P2BOMB3TIME
 288 => b"00000_0000_01_000000000000", -- load, gr0
 289 => b"00000_0000_00_000000000000", -- 0
 290 => b"00011_0000_00_001101011001", -- sub, gr0, P2BOMB3TIME
 291 => b"00110_0000_01_000000000000", -- beq
 292 => b"00000_0000_00_000110000001", -- P2EXPLOSION3INIT
 293 => b"00100_0000_01_000000000000", -- jump
 294 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 295 => b"00000_0000_01_000000000000", -- load, gr0
 296 => b"00000_0000_00_000000000000", -- 0
 297 => b"00001_0000_10_001100111100", -- store, gr0, P1BOMB1ACTIVE
 298 => b"00000_0000_00_001100111010", -- load, gr0, P1BOMB1POS
 299 => b"00001_0000_10_001100111111", -- store, gr0, P1EXPLOSION1POS
 300 => b"00000_0000_01_000000000000", -- load, gr0
 301 => b"00000_0000_00_000000000001", -- 1
 302 => b"00001_0000_10_001100111110", -- store, gr0, P1EXPLOSION1ACTIVE
 303 => b"00000_0000_01_000000000000", -- load, gr0
 304 => b"00000_0000_00_000000000010", -- 2
 305 => b"00001_0000_10_001100111101", -- store, gr0, P1EXPLOSION1TIME
 306 => b"00000_0000_00_001101011110", -- load, gr0, P1BOMBCOUNT
 307 => b"00011_0000_01_000000000000", -- sub, gr0
 308 => b"00000_0000_00_000000000001", -- 1
 309 => b"00001_0000_10_001101011110", -- store, gr0, P1BOMBCOUNT
 310 => b"00000_0100_00_001100111010", -- load, gr4, P1BOMB1POS
 311 => b"00100_0000_01_000000000000", -- jump
 312 => b"00000_0000_00_000110010011", -- EXPLODE
 313 => b"00000_0000_01_000000000000", -- load, gr0
 314 => b"00000_0000_00_000000000000", -- 0
 315 => b"00001_0000_10_001101000010", -- store, gr0, P1BOMB2ACTIVE
 316 => b"00000_0000_00_001101000000", -- load, gr0, P1BOMB2POS
 317 => b"00001_0000_10_001101000101", -- store, gr0, P1EXPLOSION2POS
 318 => b"00000_0000_01_000000000000", -- load, gr0
 319 => b"00000_0000_00_000000000001", -- 1
 320 => b"00001_0000_10_001101000100", -- store, gr0, P1EXPLOSION2ACTIVE
 321 => b"00000_0000_01_000000000000", -- load, gr0
 322 => b"00000_0000_00_000000000010", -- 2
 323 => b"00001_0000_10_001101000011", -- store, gr0, P1EXPLOSION2TIME
 324 => b"00000_0000_00_001101011110", -- load, gr0, P1BOMBCOUNT
 325 => b"00011_0000_01_000000000000", -- sub, gr0
 326 => b"00000_0000_00_000000000001", -- 1
 327 => b"00001_0000_10_001101011110", -- store, gr0, P1BOMBCOUNT
 328 => b"00000_0100_00_001101000000", -- load, gr4, P1BOMB2POS
 329 => b"00100_0000_01_000000000000", -- jump
 330 => b"00000_0000_00_000110010011", -- EXPLODE
 331 => b"00000_0000_01_000000000000", -- load, gr0
 332 => b"00000_0000_00_000000000000", -- 0
 333 => b"00001_0000_10_001101001000", -- store, gr0, P1BOMB3ACTIVE
 334 => b"00000_0000_00_001101000110", -- load, gr0, P1BOMB3POS
 335 => b"00001_0000_10_001101001011", -- store, gr0, P1EXPLOSION3POS
 336 => b"00000_0000_01_000000000000", -- load, gr0
 337 => b"00000_0000_00_000000000001", -- 1
 338 => b"00001_0000_10_001101001010", -- store, gr0, P1EXPLOSION3ACTIVE
 339 => b"00000_0000_01_000000000000", -- load, gr0
 340 => b"00000_0000_00_000000000010", -- 2
 341 => b"00001_0000_10_001101001001", -- store, gr0, P1EXPLOSION3TIME
 342 => b"00000_0000_00_001101011110", -- load, gr0, P1BOMBCOUNT
 343 => b"00011_0000_01_000000000000", -- sub, gr0
 344 => b"00000_0000_00_000000000001", -- 1
 345 => b"00001_0000_10_001101011110", -- store, gr0, P1BOMBCOUNT
 346 => b"00000_0100_00_001101000110", -- load, gr4, P1BOMB3POS
 347 => b"00100_0000_01_000000000000", -- jump
 348 => b"00000_0000_00_000110010011", -- EXPLODE
 349 => b"00000_0000_01_000000000000", -- load, gr0
 350 => b"00000_0000_00_000000000000", -- 0
 351 => b"00001_0000_10_001101001110", -- store, gr0, P2BOMB1ACTIVE
 352 => b"00000_0000_00_001101001100", -- load, gr0, P2BOMB1POS
 353 => b"00001_0000_10_001101010001", -- store, gr0, P2EXPLOSION1POS
 354 => b"00000_0000_01_000000000000", -- load, gr0
 355 => b"00000_0000_00_000000000001", -- 1
 356 => b"00001_0000_10_001101010000", -- store, gr0, P2EXPLOSION1ACTIVE
 357 => b"00000_0000_01_000000000000", -- load, gr0
 358 => b"00000_0000_00_000000000010", -- 2
 359 => b"00001_0000_10_001101001111", -- store, gr0, P2EXPLOSION1TIME
 360 => b"00000_0000_00_001101011111", -- load, gr0, P2BOMBCOUNT
 361 => b"00011_0000_01_000000000000", -- sub, gr0
 362 => b"00000_0000_00_000000000001", -- 1
 363 => b"00001_0000_10_001101011111", -- store, gr0, P2BOMBCOUNT
 364 => b"00000_0100_00_001101001100", -- load, gr4, P2BOMB1POS
 365 => b"00100_0000_01_000000000000", -- jump
 366 => b"00000_0000_00_000110010011", -- EXPLODE
 367 => b"00000_0000_01_000000000000", -- load, gr0
 368 => b"00000_0000_00_000000000000", -- 0
 369 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMB2ACTIVE
 370 => b"00000_0000_00_001101010010", -- load, gr0, P2BOMB2POS
 371 => b"00001_0000_10_001101010111", -- store, gr0, P2EXPLOSION2POS
 372 => b"00000_0000_01_000000000000", -- load, gr0
 373 => b"00000_0000_00_000000000001", -- 1
 374 => b"00001_0000_10_001101010110", -- store, gr0, P2EXPLOSION2ACTIVE
 375 => b"00000_0000_01_000000000000", -- load, gr0
 376 => b"00000_0000_00_000000000010", -- 2
 377 => b"00001_0000_10_001101010101", -- store, gr0, P2EXPLOSION2TIME
 378 => b"00000_0000_00_001101011111", -- load, gr0, P2BOMBCOUNT
 379 => b"00011_0000_01_000000000000", -- sub, gr0
 380 => b"00000_0000_00_000000000001", -- 1
 381 => b"00001_0000_10_001101011111", -- store, gr0, P2BOMBCOUNT
 382 => b"00000_0100_00_001101010010", -- load, gr4, P2BOMB2POS
 383 => b"00100_0000_01_000000000000", -- jump
 384 => b"00000_0000_00_000110010011", -- EXPLODE
 385 => b"00000_0000_01_000000000000", -- load, gr0
 386 => b"00000_0000_00_000000000000", -- 0
 387 => b"00001_0000_10_001101011010", -- store, gr0, P2BOMB3ACTIVE
 388 => b"00000_0000_00_001101011000", -- load, gr0, P2BOMB3POS
 389 => b"00001_0000_10_001101011101", -- store, gr0, P2EXPLOSION3POS
 390 => b"00000_0000_01_000000000000", -- load, gr0
 391 => b"00000_0000_00_000000000001", -- 1
 392 => b"00001_0000_10_001101011100", -- store, gr0, P2EXPLOSION3ACTIVE
 393 => b"00000_0000_01_000000000000", -- load, gr0
 394 => b"00000_0000_00_000000000010", -- 2
 395 => b"00001_0000_10_001101011011", -- store, gr0, P2EXPLOSION3TIME
 396 => b"00000_0000_00_001101011111", -- load, gr0, P2BOMBCOUNT
 397 => b"00011_0000_01_000000000000", -- sub, gr0
 398 => b"00000_0000_00_000000000001", -- 1
 399 => b"00001_0000_10_001101011111", -- store, gr0, P2BOMBCOUNT
 400 => b"00000_0100_00_001101011000", -- load, gr4, P2BOMB3POS
 401 => b"00100_0000_01_000000000000", -- jump
 402 => b"00000_0000_00_000110010011", -- EXPLODE
 403 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 404 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 405 => b"00000_0011_00_001101101011", -- load, gr3, EXPLOSION
 406 => b"10000_0010_00_000000000000", -- tpoint, gr2
 407 => b"01110_0011_00_000000000000", -- twrite, gr3
 408 => b"00010_0010_01_000000000000", -- add, gr2
 409 => b"00000_0000_00_000000000001", -- 1
 410 => b"10000_0010_00_000000000000", -- tpoint, gr2
 411 => b"01111_0000_00_000000000000", -- tread, gr0
 412 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 413 => b"00110_0000_01_000000000000", -- beq
 414 => b"00000_0000_00_000110101000", -- EXPLODELEFT
 415 => b"01110_0011_00_000000000000", -- twrite, gr3
 416 => b"00010_0010_01_000000000000", -- add, gr2
 417 => b"00000_0000_00_000000000001", -- 1
 418 => b"10000_0010_00_000000000000", -- tpoint, gr2
 419 => b"01111_0000_00_000000000000", -- tread, gr0
 420 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 421 => b"00110_0000_01_000000000000", -- beq
 422 => b"00000_0000_00_000110101000", -- EXPLODELEFT
 423 => b"01110_0011_00_000000000000", -- twrite, gr3
 424 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 425 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 426 => b"00011_0010_01_000000000000", -- sub, gr2
 427 => b"00000_0000_00_000000000001", -- 1
 428 => b"10000_0010_00_000000000000", -- tpoint, gr2
 429 => b"01111_0000_00_000000000000", -- tread, gr0
 430 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 431 => b"00110_0000_01_000000000000", -- beq
 432 => b"00000_0000_00_000110111010", -- EXPLODEDOWN
 433 => b"01110_0011_00_000000000000", -- twrite, gr3
 434 => b"00011_0010_01_000000000000", -- sub, gr2
 435 => b"00000_0000_00_000000000001", -- 1
 436 => b"10000_0010_00_000000000000", -- tpoint, gr2
 437 => b"01111_0000_00_000000000000", -- tread, gr0
 438 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 439 => b"00110_0000_01_000000000000", -- beq
 440 => b"00000_0000_00_000110111010", -- EXPLODEDOWN
 441 => b"01110_0011_00_000000000000", -- twrite, gr3
 442 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 443 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 444 => b"00010_0010_01_000000000000", -- add, gr2
 445 => b"00000_0000_00_000000001111", -- 15
 446 => b"10000_0010_00_000000000000", -- tpoint, gr2
 447 => b"01111_0000_00_000000000000", -- tread, gr0
 448 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 449 => b"00110_0000_01_000000000000", -- beq
 450 => b"00000_0000_00_000111001100", -- EXPLODEUP
 451 => b"01110_0011_00_000000000000", -- twrite, gr3
 452 => b"00010_0010_01_000000000000", -- add, gr2
 453 => b"00000_0000_00_000000001111", -- 15
 454 => b"10000_0010_00_000000000000", -- tpoint, gr2
 455 => b"01111_0000_00_000000000000", -- tread, gr0
 456 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 457 => b"00110_0000_01_000000000000", -- beq
 458 => b"00000_0000_00_000111001100", -- EXPLODEUP
 459 => b"01110_0011_00_000000000000", -- twrite, gr3
 460 => b"00001_0100_10_001101100101", -- store, gr4, MOVE
 461 => b"00000_0010_00_001101100101", -- load, gr2, MOVE
 462 => b"00011_0010_01_000000000000", -- sub, gr2
 463 => b"00000_0000_00_000000001111", -- 15
 464 => b"10000_0010_00_000000000000", -- tpoint, gr2
 465 => b"01111_0000_00_000000000000", -- tread, gr0
 466 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 467 => b"00110_0000_01_000000000000", -- beq
 468 => b"00000_0000_00_000011010001", -- TICKBOMBS
 469 => b"01110_0011_00_000000000000", -- twrite, gr3
 470 => b"00011_0010_01_000000000000", -- sub, gr2
 471 => b"00000_0000_00_000000001111", -- 15
 472 => b"10000_0010_00_000000000000", -- tpoint, gr2
 473 => b"01111_0000_00_000000000000", -- tread, gr0
 474 => b"00011_0000_00_001101101001", -- sub, gr0, WALL
 475 => b"00110_0000_01_000000000000", -- beq
 476 => b"00000_0000_00_000011010001", -- TICKBOMBS
 477 => b"01110_0011_00_000000000000", -- twrite, gr3
 478 => b"00100_0000_01_000000000000", -- jump
 479 => b"00000_0000_00_000011010001", -- TICKBOMBS
 480 => b"10101_0000_01_000000000000", -- btn1
 481 => b"00000_0000_00_000111100110", -- BTN1
 482 => b"11010_0000_01_000000000000", -- btn2
 483 => b"00000_0000_00_001001000010", -- BTN2
 484 => b"00100_0000_01_000000000000", -- jump
 485 => b"00000_0000_00_000000000100", -- BUTTON_R
 486 => b"00000_0000_00_001101011110", -- load, gr0, P1BOMBCOUNT
 487 => b"00011_0000_00_001101100000", -- sub, gr0, MAXBOMBS
 488 => b"00110_0000_01_000000000000", -- beq
 489 => b"00000_0000_00_000111100010", -- BTN1_R
 490 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 491 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 492 => b"00000_0000_00_001101100010", -- load, gr0, YPOS1
 493 => b"01000_0000_01_000000000000", -- mul, gr0
 494 => b"00000_0000_00_000000001111", -- 15
 495 => b"00010_0000_00_001101100001", -- add, gr0, XPOS1
 496 => b"10000_0000_00_000000000000", -- tpoint, gr0
 497 => b"01111_0001_00_000000000000", -- tread, gr1
 498 => b"00011_0001_00_001101101100", -- sub, gr1, EGG
 499 => b"00110_0000_01_000000000000", -- beq
 500 => b"00000_0000_00_000111100010", -- BTN1_R
 501 => b"00000_0000_00_001100111100", -- load, gr0, P1BOMB1ACTIVE
 502 => b"00011_0000_01_000000000000", -- sub, gr0
 503 => b"00000_0000_00_000000000000", -- 0
 504 => b"00110_0000_01_000000000000", -- beq
 505 => b"00000_0000_00_001000001100", -- P1PLACEBOMB1
 506 => b"00000_0000_00_001101000010", -- load, gr0, P1BOMB2ACTIVE
 507 => b"00011_0000_01_000000000000", -- sub, gr0
 508 => b"00000_0000_00_000000000000", -- 0
 509 => b"00110_0000_01_000000000000", -- beq
 510 => b"00000_0000_00_001000011110", -- P1PLACEBOMB2
 511 => b"00000_0000_00_001101001000", -- load, gr0, P1BOMB3ACTIVE
 512 => b"00011_0000_01_000000000000", -- sub, gr0
 513 => b"00000_0000_00_000000000000", -- 0
 514 => b"00110_0000_01_000000000000", -- beq
 515 => b"00000_0000_00_001000110000", -- P1PLACEBOMB3
 516 => b"00100_0000_01_000000000000", -- jump
 517 => b"00000_0000_00_000111100010", -- BTN1_R
 518 => b"00000_0000_00_001101011110", -- load, gr0, P1BOMBCOUNT
 519 => b"00010_0000_01_000000000000", -- add, gr0
 520 => b"00000_0000_00_000000000001", -- 1
 521 => b"00001_0000_10_001101011110", -- store, gr0, P1BOMBCOUNT
 522 => b"00100_0000_01_000000000000", -- jump
 523 => b"00000_0000_00_000111100010", -- BTN1_R
 524 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 525 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 526 => b"00000_0011_00_001101100010", -- load, gr3, YPOS1
 527 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 528 => b"01000_0011_01_000000000000", -- mul, gr3
 529 => b"00000_0000_00_000000001111", -- 15
 530 => b"00010_0011_00_001101100001", -- add, gr3, XPOS1
 531 => b"10000_0011_00_000000000000", -- tpoint, gr3
 532 => b"01110_0010_00_000000000000", -- twrite, gr2
 533 => b"00000_0000_01_000000000000", -- load, gr0
 534 => b"00000_0000_00_000000000001", -- 1
 535 => b"00001_0000_10_001100111100", -- store, gr0, P1BOMB1ACTIVE
 536 => b"00001_0011_10_001100111010", -- store, gr3, P1BOMB1POS
 537 => b"00000_0000_01_000000000000", -- load, gr0
 538 => b"00000_0000_00_000000010000", -- 16
 539 => b"00001_0000_10_001100111011", -- store, gr0, P1BOMB1TIME
 540 => b"00100_0000_01_000000000000", -- jump
 541 => b"00000_0000_00_001000000110", -- P1INCREASEBOMBCOUNTER
 542 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 543 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 544 => b"00000_0011_00_001101100010", -- load, gr3, YPOS1
 545 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 546 => b"01000_0011_01_000000000000", -- mul, gr3
 547 => b"00000_0000_00_000000001111", -- 15
 548 => b"00010_0011_00_001101100001", -- add, gr3, XPOS1
 549 => b"10000_0011_00_000000000000", -- tpoint, gr3
 550 => b"01110_0010_00_000000000000", -- twrite, gr2
 551 => b"00000_0000_01_000000000000", -- load, gr0
 552 => b"00000_0000_00_000000000001", -- 1
 553 => b"00001_0000_10_001101000010", -- store, gr0, P1BOMB2ACTIVE
 554 => b"00001_0011_10_001101000000", -- store, gr3, P1BOMB2POS
 555 => b"00000_0000_01_000000000000", -- load, gr0
 556 => b"00000_0000_00_000000010000", -- 16
 557 => b"00001_0000_10_001101000001", -- store, gr0, P1BOMB2TIME
 558 => b"00100_0000_01_000000000000", -- jump
 559 => b"00000_0000_00_001000000110", -- P1INCREASEBOMBCOUNTER
 560 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 561 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 562 => b"00000_0011_00_001101100010", -- load, gr3, YPOS1
 563 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 564 => b"01000_0011_01_000000000000", -- mul, gr3
 565 => b"00000_0000_00_000000001111", -- 15
 566 => b"00010_0011_00_001101100001", -- add, gr3, XPOS1
 567 => b"10000_0011_00_000000000000", -- tpoint, gr3
 568 => b"01110_0010_00_000000000000", -- twrite, gr2
 569 => b"00000_0000_01_000000000000", -- load, gr0
 570 => b"00000_0000_00_000000000001", -- 1
 571 => b"00001_0000_10_001101001000", -- store, gr0, P1BOMB3ACTIVE
 572 => b"00001_0011_10_001101000110", -- store, gr3, P1BOMB3POS
 573 => b"00000_0000_01_000000000000", -- load, gr0
 574 => b"00000_0000_00_000000010000", -- 16
 575 => b"00001_0000_10_001101000111", -- store, gr0, P1BOMB3TIME
 576 => b"00100_0000_01_000000000000", -- jump
 577 => b"00000_0000_00_001000000110", -- P1INCREASEBOMBCOUNTER
 578 => b"00000_0000_00_001101011111", -- load, gr0, P2BOMBCOUNT
 579 => b"00011_0000_00_001101100000", -- sub, gr0, MAXBOMBS
 580 => b"00110_0000_01_000000000000", -- beq
 581 => b"00000_0000_00_000111100100", -- BTN2_R
 582 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 583 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 584 => b"00000_0000_00_001101100100", -- load, gr0, YPOS2
 585 => b"01000_0000_01_000000000000", -- mul, gr0
 586 => b"00000_0000_00_000000001111", -- 15
 587 => b"00010_0000_00_001101100011", -- add, gr0, XPOS2
 588 => b"10000_0000_00_000000000000", -- tpoint, gr0
 589 => b"01111_0001_00_000000000000", -- tread, gr1
 590 => b"00011_0001_00_001101101100", -- sub, gr1, EGG
 591 => b"00110_0000_01_000000000000", -- beq
 592 => b"00000_0000_00_000111100100", -- BTN2_R
 593 => b"00000_0000_00_001101001110", -- load, gr0, P2BOMB1ACTIVE
 594 => b"00011_0000_01_000000000000", -- sub, gr0
 595 => b"00000_0000_00_000000000000", -- 0
 596 => b"00110_0000_01_000000000000", -- beq
 597 => b"00000_0000_00_001001100110", -- P2PLACEBOMB1
 598 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMB2ACTIVE
 599 => b"00011_0000_01_000000000000", -- sub, gr0
 600 => b"00000_0000_00_000000000000", -- 0
 601 => b"00110_0000_01_000000000000", -- beq
 602 => b"00000_0000_00_001001111000", -- P2PLACEBOMB2
 603 => b"00000_0000_00_001101011010", -- load, gr0, P2BOMB3ACTIVE
 604 => b"00011_0000_01_000000000000", -- sub, gr0
 605 => b"00000_0000_00_000000000000", -- 0
 606 => b"00110_0000_01_000000000000", -- beq
 607 => b"00000_0000_00_001010001010", -- P2PLACEBOMB3
 608 => b"00000_0000_00_001101011111", -- load, gr0, P2BOMBCOUNT
 609 => b"00010_0000_01_000000000000", -- add, gr0
 610 => b"00000_0000_00_000000000001", -- 1
 611 => b"00001_0000_10_001101011111", -- store, gr0, P2BOMBCOUNT
 612 => b"00100_0000_01_000000000000", -- jump
 613 => b"00000_0000_00_000111100100", -- BTN2_R
 614 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 615 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 616 => b"00000_0011_00_001101100100", -- load, gr3, YPOS2
 617 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 618 => b"01000_0011_01_000000000000", -- mul, gr3
 619 => b"00000_0000_00_000000001111", -- 15
 620 => b"00010_0011_00_001101100011", -- add, gr3, XPOS2
 621 => b"10000_0011_00_000000000000", -- tpoint, gr3
 622 => b"01110_0010_00_000000000000", -- twrite, gr2
 623 => b"00000_0000_01_000000000000", -- load, gr0
 624 => b"00000_0000_00_000000000001", -- 1
 625 => b"00001_0000_10_001101001110", -- store, gr0, P2BOMB1ACTIVE
 626 => b"00001_0011_10_001101001100", -- store, gr3, P2BOMB1POS
 627 => b"00000_0000_01_000000000000", -- load, gr0
 628 => b"00000_0000_00_000000010000", -- 16
 629 => b"00001_0000_10_001101001101", -- store, gr0, P2BOMB1TIME
 630 => b"00100_0000_01_000000000000", -- jump
 631 => b"00000_0000_00_001001100000", -- P2INCREASEBOMBCOUNTER
 632 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 633 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 634 => b"00000_0011_00_001101100100", -- load, gr3, YPOS2
 635 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 636 => b"01000_0011_01_000000000000", -- mul, gr3
 637 => b"00000_0000_00_000000001111", -- 15
 638 => b"00010_0011_00_001101100011", -- add, gr3, XPOS2
 639 => b"10000_0011_00_000000000000", -- tpoint, gr3
 640 => b"01110_0010_00_000000000000", -- twrite, gr2
 641 => b"00000_0000_01_000000000000", -- load, gr0
 642 => b"00000_0000_00_000000000001", -- 1
 643 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMB2ACTIVE
 644 => b"00001_0011_10_001101010010", -- store, gr3, P2BOMB2POS
 645 => b"00000_0000_01_000000000000", -- load, gr0
 646 => b"00000_0000_00_000000010000", -- 16
 647 => b"00001_0000_10_001101010011", -- store, gr0, P2BOMB2TIME
 648 => b"00100_0000_01_000000000000", -- jump
 649 => b"00000_0000_00_001001100000", -- P2INCREASEBOMBCOUNTER
 650 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 651 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 652 => b"00000_0011_00_001101100100", -- load, gr3, YPOS2
 653 => b"00000_0010_00_001101101100", -- load, gr2, EGG
 654 => b"01000_0011_01_000000000000", -- mul, gr3
 655 => b"00000_0000_00_000000001111", -- 15
 656 => b"00010_0011_00_001101100011", -- add, gr3, XPOS2
 657 => b"10000_0011_00_000000000000", -- tpoint, gr3
 658 => b"01110_0010_00_000000000000", -- twrite, gr2
 659 => b"00000_0000_01_000000000000", -- load, gr0
 660 => b"00000_0000_00_000000000001", -- 1
 661 => b"00001_0000_10_001101011010", -- store, gr0, P2BOMB3ACTIVE
 662 => b"00001_0011_10_001101011000", -- store, gr3, P2BOMB3POS
 663 => b"00000_0000_01_000000000000", -- load, gr0
 664 => b"00000_0000_00_000000010000", -- 16
 665 => b"00001_0000_10_001101011001", -- store, gr0, P2BOMB3TIME
 666 => b"00100_0000_01_000000000000", -- jump
 667 => b"00000_0000_00_001001100000", -- P2INCREASEBOMBCOUNTER
 668 => b"00100_0000_01_000000000000", -- jump
 669 => b"00000_0000_00_001100111000", -- COUNT1
 670 => b"10001_0000_01_000000000000", -- joy1r
 671 => b"00000_0000_00_001010110000", -- P1R
 672 => b"10011_0000_01_000000000000", -- joy1l
 673 => b"00000_0000_00_001011010010", -- P1L
 674 => b"10010_0000_01_000000000000", -- joy1u
 675 => b"00000_0000_00_001011000001", -- P1U
 676 => b"10100_0000_01_000000000000", -- joy1d
 677 => b"00000_0000_00_001011100011", -- P1D
 678 => b"10110_0000_01_000000000000", -- joy2r
 679 => b"00000_0000_00_001011110100", -- P2R
 680 => b"11000_0000_01_000000000000", -- joy2l
 681 => b"00000_0000_00_001100010110", -- P2L
 682 => b"10111_0000_01_000000000000", -- joy2u
 683 => b"00000_0000_00_001100000101", -- P2U
 684 => b"11001_0000_01_000000000000", -- joy2d
 685 => b"00000_0000_00_001100100111", -- P2D
 686 => b"00100_0000_01_000000000000", -- jump
 687 => b"00000_0000_00_000000000010", -- CONTROL_R
 688 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 689 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 690 => b"00000_0000_00_001101100010", -- load, gr0, YPOS1
 691 => b"01000_0000_01_000000000000", -- mul, gr0
 692 => b"00000_0000_00_000000001111", -- 15
 693 => b"00010_0000_00_001101100001", -- add, gr0, XPOS1
 694 => b"00010_0000_01_000000000000", -- add, gr0
 695 => b"00000_0000_00_000000000001", -- 1
 696 => b"10000_0000_00_000000000000", -- tpoint, gr0
 697 => b"01111_0001_00_000000000000", -- tread, gr1
 698 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 699 => b"00111_0000_01_000000000000", -- bne
 700 => b"00000_0000_00_001010100010", -- J1
 701 => b"00010_1100_01_000000000000", -- add, gr12
 702 => b"00000_0000_00_000000000001", -- 1
 703 => b"00100_0000_01_000000000000", -- jump
 704 => b"00000_0000_00_001010100010", -- J1
 705 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 706 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 707 => b"00000_0000_00_001101100010", -- load, gr0, YPOS1
 708 => b"00011_0000_01_000000000000", -- sub, gr0
 709 => b"00000_0000_00_000000000001", -- 1
 710 => b"01000_0000_01_000000000000", -- mul, gr0
 711 => b"00000_0000_00_000000001111", -- 15
 712 => b"00010_0000_00_001101100001", -- add, gr0, XPOS1
 713 => b"10000_0000_00_000000000000", -- tpoint, gr0
 714 => b"01111_0001_00_000000000000", -- tread, gr1
 715 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 716 => b"00111_0000_01_000000000000", -- bne
 717 => b"00000_0000_00_001010100110", -- J2
 718 => b"00011_1101_01_000000000000", -- sub, gr13
 719 => b"00000_0000_00_000000000001", -- 1
 720 => b"00100_0000_01_000000000000", -- jump
 721 => b"00000_0000_00_001010100110", -- J2
 722 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 723 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 724 => b"00000_0000_00_001101100010", -- load, gr0, YPOS1
 725 => b"01000_0000_01_000000000000", -- mul, gr0
 726 => b"00000_0000_00_000000001111", -- 15
 727 => b"00010_0000_00_001101100001", -- add, gr0, XPOS1
 728 => b"00011_0000_01_000000000000", -- sub, gr0
 729 => b"00000_0000_00_000000000001", -- 1
 730 => b"10000_0000_00_000000000000", -- tpoint, gr0
 731 => b"01111_0001_00_000000000000", -- tread, gr1
 732 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 733 => b"00111_0000_01_000000000000", -- bne
 734 => b"00000_0000_00_001010100010", -- J1
 735 => b"00011_1100_01_000000000000", -- sub, gr12
 736 => b"00000_0000_00_000000000001", -- 1
 737 => b"00100_0000_01_000000000000", -- jump
 738 => b"00000_0000_00_001010100010", -- J1
 739 => b"00001_1100_10_001101100001", -- store, gr12, XPOS1
 740 => b"00001_1101_10_001101100010", -- store, gr13, YPOS1
 741 => b"00000_0000_00_001101100010", -- load, gr0, YPOS1
 742 => b"00010_0000_01_000000000000", -- add, gr0
 743 => b"00000_0000_00_000000000001", -- 1
 744 => b"01000_0000_01_000000000000", -- mul, gr0
 745 => b"00000_0000_00_000000001111", -- 15
 746 => b"00010_0000_00_001101100001", -- add, gr0, XPOS1
 747 => b"10000_0000_00_000000000000", -- tpoint, gr0
 748 => b"01111_0001_00_000000000000", -- tread, gr1
 749 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 750 => b"00111_0000_01_000000000000", -- bne
 751 => b"00000_0000_00_001010100110", -- J2
 752 => b"00010_1101_01_000000000000", -- add, gr13
 753 => b"00000_0000_00_000000000001", -- 1
 754 => b"00100_0000_01_000000000000", -- jump
 755 => b"00000_0000_00_001010100110", -- J2
 756 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 757 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 758 => b"00000_0000_00_001101100100", -- load, gr0, YPOS2
 759 => b"01000_0000_01_000000000000", -- mul, gr0
 760 => b"00000_0000_00_000000001111", -- 15
 761 => b"00010_0000_00_001101100011", -- add, gr0, XPOS2
 762 => b"00010_0000_01_000000000000", -- add, gr0
 763 => b"00000_0000_00_000000000001", -- 1
 764 => b"10000_0000_00_000000000000", -- tpoint, gr0
 765 => b"01111_0001_00_000000000000", -- tread, gr1
 766 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 767 => b"00111_0000_01_000000000000", -- bne
 768 => b"00000_0000_00_001010101010", -- J3
 769 => b"00010_1110_01_000000000000", -- add, gr14
 770 => b"00000_0000_00_000000000001", -- 1
 771 => b"00100_0000_01_000000000000", -- jump
 772 => b"00000_0000_00_001010101010", -- J3
 773 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 774 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 775 => b"00000_0000_00_001101100100", -- load, gr0, YPOS2
 776 => b"00011_0000_01_000000000000", -- sub, gr0
 777 => b"00000_0000_00_000000000001", -- 1
 778 => b"01000_0000_01_000000000000", -- mul, gr0
 779 => b"00000_0000_00_000000001111", -- 15
 780 => b"00010_0000_00_001101100011", -- add, gr0, XPOS2
 781 => b"10000_0000_00_000000000000", -- tpoint, gr0
 782 => b"01111_0001_00_000000000000", -- tread, gr1
 783 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 784 => b"00111_0000_01_000000000000", -- bne
 785 => b"00000_0000_00_000000000010", -- CONTROL_R
 786 => b"00011_1111_01_000000000000", -- sub, gr15
 787 => b"00000_0000_00_000000000001", -- 1
 788 => b"00100_0000_01_000000000000", -- jump
 789 => b"00000_0000_00_000000000010", -- CONTROL_R
 790 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 791 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 792 => b"00000_0000_00_001101100100", -- load, gr0, YPOS2
 793 => b"01000_0000_01_000000000000", -- mul, gr0
 794 => b"00000_0000_00_000000001111", -- 15
 795 => b"00010_0000_00_001101100011", -- add, gr0, XPOS2
 796 => b"00011_0000_01_000000000000", -- sub, gr0
 797 => b"00000_0000_00_000000000001", -- 1
 798 => b"10000_0000_00_000000000000", -- tpoint, gr0
 799 => b"01111_0001_00_000000000000", -- tread, gr1
 800 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 801 => b"00111_0000_01_000000000000", -- bne
 802 => b"00000_0000_00_001010101010", -- J3
 803 => b"00011_1110_01_000000000000", -- sub, gr14
 804 => b"00000_0000_00_000000000001", -- 1
 805 => b"00100_0000_01_000000000000", -- jump
 806 => b"00000_0000_00_001010101010", -- J3
 807 => b"00001_1110_10_001101100011", -- store, gr14, XPOS2
 808 => b"00001_1111_10_001101100100", -- store, gr15, YPOS2
 809 => b"00000_0000_00_001101100100", -- load, gr0, YPOS2
 810 => b"00010_0000_01_000000000000", -- add, gr0
 811 => b"00000_0000_00_000000000001", -- 1
 812 => b"01000_0000_01_000000000000", -- mul, gr0
 813 => b"00000_0000_00_000000001111", -- 15
 814 => b"00010_0000_00_001101100011", -- add, gr0, XPOS2
 815 => b"10000_0000_00_000000000000", -- tpoint, gr0
 816 => b"01111_0001_00_000000000000", -- tread, gr1
 817 => b"00011_0001_00_001101101000", -- sub, gr1, GRASS
 818 => b"00111_0000_01_000000000000", -- bne
 819 => b"00000_0000_00_000000000010", -- CONTROL_R
 820 => b"00010_1111_01_000000000000", -- add, gr15
 821 => b"00000_0000_00_000000000001", -- 1
 822 => b"00100_0000_01_000000000000", -- jump
 823 => b"00000_0000_00_000000000010", -- CONTROL_R
 824 => b"00100_0000_01_000000000000", -- jump
 825 => b"00000_0000_00_001010011110", -- COUNT_R
 826 => b"00000_0000_00_000000000000", -- 0
 827 => b"00000_0000_00_000000000000", -- 0
 828 => b"00000_0000_00_000000000000", -- 0
 829 => b"00000_0000_00_000000000000", -- 0
 830 => b"00000_0000_00_000000000000", -- 0
 831 => b"00000_0000_00_000000000000", -- 0
 832 => b"00000_0000_00_000000000000", -- 0
 833 => b"00000_0000_00_000000000000", -- 0
 834 => b"00000_0000_00_000000000000", -- 0
 835 => b"00000_0000_00_000000000000", -- 0
 836 => b"00000_0000_00_000000000000", -- 0
 837 => b"00000_0000_00_000000000000", -- 0
 838 => b"00000_0000_00_000000000000", -- 0
 839 => b"00000_0000_00_000000000000", -- 0
 840 => b"00000_0000_00_000000000000", -- 0
 841 => b"00000_0000_00_000000000000", -- 0
 842 => b"00000_0000_00_000000000000", -- 0
 843 => b"00000_0000_00_000000000000", -- 0
 844 => b"00000_0000_00_000000000000", -- 0
 845 => b"00000_0000_00_000000000000", -- 0
 846 => b"00000_0000_00_000000000000", -- 0
 847 => b"00000_0000_00_000000000000", -- 0
 848 => b"00000_0000_00_000000000000", -- 0
 849 => b"00000_0000_00_000000000000", -- 0
 850 => b"00000_0000_00_000000000000", -- 0
 851 => b"00000_0000_00_000000000000", -- 0
 852 => b"00000_0000_00_000000000000", -- 0
 853 => b"00000_0000_00_000000000000", -- 0
 854 => b"00000_0000_00_000000000000", -- 0
 855 => b"00000_0000_00_000000000000", -- 0
 856 => b"00000_0000_00_000000000000", -- 0
 857 => b"00000_0000_00_000000000000", -- 0
 858 => b"00000_0000_00_000000000000", -- 0
 859 => b"00000_0000_00_000000000000", -- 0
 860 => b"00000_0000_00_000000000000", -- 0
 861 => b"00000_0000_00_000000000000", -- 0
 862 => b"00000_0000_00_000000000000", -- 0
 863 => b"00000_0000_00_000000000000", -- 0
 864 => b"00000_0000_00_000000000011", -- 3
 865 => b"00000_0000_00_000000000000", -- 0
 866 => b"00000_0000_00_000000000000", -- 0
 867 => b"00000_0000_00_000000000000", -- 0
 868 => b"00000_0000_00_000000000000", -- 0
 869 => b"00000_0000_00_000000000000", -- 0
 870 => b"00000_0000_00_000000000000", -- 0
 871 => b"00000_0000_00_000000000000", -- 0
 872 => b"00000_0000_00_000000000000", -- 0
 873 => b"00000_0000_00_000000000001", -- 1
 874 => b"00000_0000_00_000000000010", -- 2
 875 => b"00000_0000_00_000000000011", -- 3
 876 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
