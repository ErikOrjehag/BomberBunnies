library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity MICRO_MEMORY is
  port (
    uAddr : in unsigned(8 downto 0);
    uData : out std_logic_vector(29 downto 0));
end MICRO_MEMORY;

architecture Behavioral of MICRO_MEMORY is

-- micro Memory
type u_mem_t is array (0 to 511) of std_logic_vector(29 downto 0);
constant u_mem_c : u_mem_t := (
  -- AR 0110
       --   ALU   TB   FB  S P LC  SEQ  uADR
    0  => b"0000_0100_0001_0_0_00_00000_000000000",  -- H�mtfas
    1  => b"0000_0011_0010_0_1_00_00000_000000000",
    
    2  => b"0000_0000_0000_0_0_00_00010_000000000",  -- Start
    
    3  => b"0000_0010_0001_0_0_00_00001_000000000",  -- Direktadressering
    
    4  => b"0000_0100_0001_0_1_00_00001_000000000",  -- Immediate
    
    5  => b"0000_0010_0001_0_0_00_00000_000000000",  -- Indirekt adressering
    6  => b"0000_0011_0001_0_0_00_00001_000000000",
    
    7  => b"0000_0110_0000_0_0_00_00000_000000000",  -- Indexerad adressering
    8  => b"1000_0101_0000_0_0_00_00000_000000000",
    9  => b"0000_0110_0001_0_0_00_00001_000000000",
    
    
    10 => b"0000_0011_0101_0_0_00_00011_000000000",  -- LOAD (GRx, M, ADDR)

    11 => b"0000_0010_0001_0_0_00_00000_000000000",  -- STORE (GRx, M, ADDR)
    12 => b"0000_0101_0011_0_0_00_00011_000000000",
    
    13 => b"0001_0011_0000_0_0_00_00000_000000000",  -- ADD (GRx, M, ADDR)
    14 => b"0100_0101_0000_0_0_00_00000_000000000",
    15 => b"0000_0110_0101_0_0_00_00011_000000000",
    
    16 => b"0001_0101_0000_0_0_00_00000_000000000",  -- SUB (GRx, M, ADDR)
    17 => b"0101_0011_0000_0_0_00_00000_000000000",
    18 => b"0000_0110_0101_0_0_00_00011_000000000",
    
    19 => b"0000_0011_0100_0_0_00_00011_000000000",  -- JUMP
    
    20 => b"0000_0011_0000_0_0_00_00000_000000000",  -- SLEEP
    21 => b"0000_0000_0000_0_0_10_00000_000000000",
    22 => b"0000_0000_0000_0_0_01_00000_000000000",
    23 => b"0000_0000_0000_0_0_00_01100_000010101",
    24 => b"0000_0000_0000_0_0_00_00011_000000000",

    25 => b"0000_0000_0000_0_0_00_01000_000010010",  -- BEQ (g�r till JUMP om 
    26 => b"0000_0000_0000_0_0_00_00011_000000000",  -- z = 1.)

    27 => b"0000_0000_0000_0_0_00_00100_000010010",  -- BNE (g�r till JUMP om 
    28 => b"0000_0000_0000_0_1_00_00011_000000000",  -- z = 0, annars PC+1.)

    -- Stort h�l h�r!

    34 => b"0000_0101_1000_0_0_00_00011_000000000",  -- GRx till tileWrite,
    --35 => b"0000_0000_0000_0_0_00_00011_000000000",

    36 => b"0000_1000_0101_0_0_00_00011_000000000",  -- tileRead to GRx
    --37 => b"0000_0000_0000_0_0_00_00011_000000000",

    38 => b"0000_0101_1001_0_0_00_00011_000000000",  -- GRx to tilePointer

    39 => b"0000_0000_0000_0_0_00_10000_000010011",  -- JOY1R (g�r till JUMP om 
    40 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j1r = 1.)

    41 => b"0000_0000_0000_0_0_00_10001_000010011",  -- JOY1U (g�r till JUMP om
    42 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j1u = 1.)

    43 => b"0000_0000_0000_0_0_00_10010_000010011",  -- JOY1L (g�r till JUMP om
    44 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j1l = 1.)

    45 => b"0000_0000_0000_0_0_00_10011_000010011",  -- JOY1D (g�r till JUMP om
    46 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j1d = 1.)

    47 => b"0000_0000_0000_0_0_00_10100_000010011",  -- BTN1 (g�r till JUMP om
    48 => b"0000_0000_0000_0_0_00_00011_000000000",  -- b1 = 1.)
    
    49 => b"0000_0000_0000_0_0_00_10101_000010011",  -- JOY2R (g�r till JUMP om
    50 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j2r = 1.)
    
    51 => b"0000_0000_0000_0_0_00_10110_000010011",  -- JOY2U (g�r till JUMP om
    52 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j2u = 1.)

    53 => b"0000_0000_0000_0_0_00_10111_000010011",  -- JOY2L (g�r till JUMP om
    54 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j2l = 1.)

    56 => b"0000_0000_0000_0_0_00_11000_000010011",  -- JOY2D (g�r till JUMP om
    57 => b"0000_0000_0000_0_0_00_00011_000000000",  -- j2d = 1.)

    58 => b"0000_0000_0000_0_0_00_11001_000010011",  -- BTN2 (g�r till JUMP om
    59 => b"0000_0000_0000_0_0_00_00011_000000000",  -- b2 = 1.)
    
    others => (others => '0')
  );

signal uMem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= uMem(to_integer(uAddr));

end Behavioral;
