library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr
0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000001001011", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000000001000", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000000010", -- MAIN
   8 => b"10101_0000_01_000000000000", -- btn1
   9 => b"00000_0000_00_000000001110", -- BTN1
  10 => b"11010_0000_01_000000000000", -- btn2
  11 => b"00000_0000_00_000000101100", -- BTN2
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000000000110", -- BUTTON_R
  14 => b"00000_0000_00_000011101001", -- load, gr0, BOMBS1
  15 => b"00011_0000_00_000011101011", -- sub, gr0, MAXBOMBS
  16 => b"00110_0000_01_000000000000", -- beq
  17 => b"00000_0000_00_000000001010", -- BTN1_R
  18 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
  19 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
  20 => b"00000_0000_00_000011110010", -- load, gr0, YPOS1
  21 => b"01000_0000_01_000000000000", -- mul, gr0
  22 => b"00000_0000_00_000000001111", -- 15
  23 => b"00010_0000_00_000011110001", -- add, gr0, XPOS1
  24 => b"10000_0000_00_000000000000", -- tpoint, gr0
  25 => b"01111_0001_00_000000000000", -- tread, gr1
  26 => b"00011_0001_00_000011110000", -- sub, gr1, EGG
  27 => b"00110_0000_01_000000000000", -- beq
  28 => b"00000_0000_00_000000001100", -- BTN2_R
  29 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
  30 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
  31 => b"00000_0011_00_000011110010", -- load, gr3, YPOS1
  32 => b"00000_0010_00_000011110000", -- load, gr2, EGG
  33 => b"01000_0011_01_000000000000", -- mul, gr3
  34 => b"00000_0000_00_000000001111", -- 15
  35 => b"00010_0011_00_000011110001", -- add, gr3, XPOS1
  36 => b"10000_0011_00_000000000000", -- tpoint, gr3
  37 => b"01110_0010_00_000000000000", -- twrite, gr2
  38 => b"00000_0000_00_000011101001", -- load, gr0, BOMBS1
  39 => b"00010_0000_01_000000000000", -- add, gr0
  40 => b"00000_0000_00_000000000001", -- 1
  41 => b"00001_0000_10_000011101001", -- store, gr0, BOMBS1
  42 => b"00100_0000_01_000000000000", -- jump
  43 => b"00000_0000_00_000000001010", -- BTN1_R
  44 => b"00000_0000_00_000011101010", -- load, gr0, BOMBS2
  45 => b"00011_0000_00_000011101011", -- sub, gr0, MAXBOMBS
  46 => b"00110_0000_01_000000000000", -- beq
  47 => b"00000_0000_00_000000001100", -- BTN2_R
  48 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
  49 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
  50 => b"00000_0000_00_000011110100", -- load, gr0, YPOS2
  51 => b"01000_0000_01_000000000000", -- mul, gr0
  52 => b"00000_0000_00_000000001111", -- 15
  53 => b"00010_0000_00_000011110011", -- add, gr0, XPOS2
  54 => b"10000_0000_00_000000000000", -- tpoint, gr0
  55 => b"01111_0001_00_000000000000", -- tread, gr1
  56 => b"00011_0001_00_000011110000", -- sub, gr1, EGG
  57 => b"00110_0000_01_000000000000", -- beq
  58 => b"00000_0000_00_000000001100", -- BTN2_R
  59 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
  60 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
  61 => b"00000_0011_00_000011110100", -- load, gr3, YPOS2
  62 => b"00000_0010_00_000011110000", -- load, gr2, EGG
  63 => b"01000_0011_01_000000000000", -- mul, gr3
  64 => b"00000_0000_00_000000001111", -- 15
  65 => b"00010_0011_00_000011110011", -- add, gr3, XPOS2
  66 => b"10000_0011_00_000000000000", -- tpoint, gr3
  67 => b"01110_0010_00_000000000000", -- twrite, gr2
  68 => b"00000_0000_00_000011101010", -- load, gr0, BOMBS2
  69 => b"00010_0000_01_000000000000", -- add, gr0
  70 => b"00000_0000_00_000000000001", -- 1
  71 => b"00001_0000_10_000011101010", -- store, gr0, BOMBS2
  72 => b"00100_0000_01_000000000000", -- jump
  73 => b"00000_0000_00_000000001100", -- BTN2_R
  74 => b"00000_0000_00_000000000000", -- 0
  75 => b"00100_0000_01_000000000000", -- jump
  76 => b"00000_0000_00_000011100111", -- COUNT1
  77 => b"10001_0000_01_000000000000", -- joy1r
  78 => b"00000_0000_00_000001011111", -- P1R
  79 => b"10011_0000_01_000000000000", -- joy1l
  80 => b"00000_0000_00_000010000001", -- P1L
  81 => b"10010_0000_01_000000000000", -- joy1u
  82 => b"00000_0000_00_000001110000", -- P1U
  83 => b"10100_0000_01_000000000000", -- joy1d
  84 => b"00000_0000_00_000010010010", -- P1D
  85 => b"10110_0000_01_000000000000", -- joy2r
  86 => b"00000_0000_00_000010100011", -- P2R
  87 => b"11000_0000_01_000000000000", -- joy2l
  88 => b"00000_0000_00_000011000101", -- P2L
  89 => b"10111_0000_01_000000000000", -- joy2u
  90 => b"00000_0000_00_000010110100", -- P2U
  91 => b"11001_0000_01_000000000000", -- joy2d
  92 => b"00000_0000_00_000011010110", -- P2D
  93 => b"00100_0000_01_000000000000", -- jump
  94 => b"00000_0000_00_000000000100", -- CONTROL_R
  95 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
  96 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
  97 => b"00000_0000_00_000011110010", -- load, gr0, YPOS1
  98 => b"01000_0000_01_000000000000", -- mul, gr0
  99 => b"00000_0000_00_000000001111", -- 15
 100 => b"00010_0000_00_000011110001", -- add, gr0, XPOS1
 101 => b"00010_0000_01_000000000000", -- add, gr0
 102 => b"00000_0000_00_000000000001", -- 1
 103 => b"10000_0000_00_000000000000", -- tpoint, gr0
 104 => b"01111_0001_00_000000000000", -- tread, gr1
 105 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 106 => b"00111_0000_01_000000000000", -- bne
 107 => b"00000_0000_00_000001010001", -- J1
 108 => b"00010_1100_01_000000000000", -- add, gr12
 109 => b"00000_0000_00_000000000001", -- 1
 110 => b"00100_0000_01_000000000000", -- jump
 111 => b"00000_0000_00_000001010001", -- J1
 112 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
 113 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
 114 => b"00000_0000_00_000011110010", -- load, gr0, YPOS1
 115 => b"00011_0000_01_000000000000", -- sub, gr0
 116 => b"00000_0000_00_000000000001", -- 1
 117 => b"01000_0000_01_000000000000", -- mul, gr0
 118 => b"00000_0000_00_000000001111", -- 15
 119 => b"00010_0000_00_000011110001", -- add, gr0, XPOS1
 120 => b"10000_0000_00_000000000000", -- tpoint, gr0
 121 => b"01111_0001_00_000000000000", -- tread, gr1
 122 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 123 => b"00111_0000_01_000000000000", -- bne
 124 => b"00000_0000_00_000001010101", -- J2
 125 => b"00011_1101_01_000000000000", -- sub, gr13
 126 => b"00000_0000_00_000000000001", -- 1
 127 => b"00100_0000_01_000000000000", -- jump
 128 => b"00000_0000_00_000001010101", -- J2
 129 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
 130 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
 131 => b"00000_0000_00_000011110010", -- load, gr0, YPOS1
 132 => b"01000_0000_01_000000000000", -- mul, gr0
 133 => b"00000_0000_00_000000001111", -- 15
 134 => b"00010_0000_00_000011110001", -- add, gr0, XPOS1
 135 => b"00011_0000_01_000000000000", -- sub, gr0
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0000_00_000000000000", -- tpoint, gr0
 138 => b"01111_0001_00_000000000000", -- tread, gr1
 139 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000001010001", -- J1
 142 => b"00011_1100_01_000000000000", -- sub, gr12
 143 => b"00000_0000_00_000000000001", -- 1
 144 => b"00100_0000_01_000000000000", -- jump
 145 => b"00000_0000_00_000001010001", -- J1
 146 => b"00001_1100_10_000011110001", -- store, gr12, XPOS1
 147 => b"00001_1101_10_000011110010", -- store, gr13, YPOS1
 148 => b"00000_0000_00_000011110010", -- load, gr0, YPOS1
 149 => b"00010_0000_01_000000000000", -- add, gr0
 150 => b"00000_0000_00_000000000001", -- 1
 151 => b"01000_0000_01_000000000000", -- mul, gr0
 152 => b"00000_0000_00_000000001111", -- 15
 153 => b"00010_0000_00_000011110001", -- add, gr0, XPOS1
 154 => b"10000_0000_00_000000000000", -- tpoint, gr0
 155 => b"01111_0001_00_000000000000", -- tread, gr1
 156 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000001010101", -- J2
 159 => b"00010_1101_01_000000000000", -- add, gr13
 160 => b"00000_0000_00_000000000001", -- 1
 161 => b"00100_0000_01_000000000000", -- jump
 162 => b"00000_0000_00_000001010101", -- J2
 163 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
 164 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
 165 => b"00000_0000_00_000011110100", -- load, gr0, YPOS2
 166 => b"01000_0000_01_000000000000", -- mul, gr0
 167 => b"00000_0000_00_000000001111", -- 15
 168 => b"00010_0000_00_000011110011", -- add, gr0, XPOS2
 169 => b"00010_0000_01_000000000000", -- add, gr0
 170 => b"00000_0000_00_000000000001", -- 1
 171 => b"10000_0000_00_000000000000", -- tpoint, gr0
 172 => b"01111_0001_00_000000000000", -- tread, gr1
 173 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000001011001", -- J3
 176 => b"00010_1110_01_000000000000", -- add, gr14
 177 => b"00000_0000_00_000000000001", -- 1
 178 => b"00100_0000_01_000000000000", -- jump
 179 => b"00000_0000_00_000001011001", -- J3
 180 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
 181 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
 182 => b"00000_0000_00_000011110100", -- load, gr0, YPOS2
 183 => b"00011_0000_01_000000000000", -- sub, gr0
 184 => b"00000_0000_00_000000000001", -- 1
 185 => b"01000_0000_01_000000000000", -- mul, gr0
 186 => b"00000_0000_00_000000001111", -- 15
 187 => b"00010_0000_00_000011110011", -- add, gr0, XPOS2
 188 => b"10000_0000_00_000000000000", -- tpoint, gr0
 189 => b"01111_0001_00_000000000000", -- tread, gr1
 190 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000000100", -- CONTROL_R
 193 => b"00011_1111_01_000000000000", -- sub, gr15
 194 => b"00000_0000_00_000000000001", -- 1
 195 => b"00100_0000_01_000000000000", -- jump
 196 => b"00000_0000_00_000000000100", -- CONTROL_R
 197 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
 198 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
 199 => b"00000_0000_00_000011110100", -- load, gr0, YPOS2
 200 => b"01000_0000_01_000000000000", -- mul, gr0
 201 => b"00000_0000_00_000000001111", -- 15
 202 => b"00010_0000_00_000011110011", -- add, gr0, XPOS2
 203 => b"00011_0000_01_000000000000", -- sub, gr0
 204 => b"00000_0000_00_000000000001", -- 1
 205 => b"10000_0000_00_000000000000", -- tpoint, gr0
 206 => b"01111_0001_00_000000000000", -- tread, gr1
 207 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 208 => b"00111_0000_01_000000000000", -- bne
 209 => b"00000_0000_00_000001011001", -- J3
 210 => b"00011_1110_01_000000000000", -- sub, gr14
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00100_0000_01_000000000000", -- jump
 213 => b"00000_0000_00_000001011001", -- J3
 214 => b"00001_1110_10_000011110011", -- store, gr14, XPOS2
 215 => b"00001_1111_10_000011110100", -- store, gr15, YPOS2
 216 => b"00000_0000_00_000011110100", -- load, gr0, YPOS2
 217 => b"00010_0000_01_000000000000", -- add, gr0
 218 => b"00000_0000_00_000000000001", -- 1
 219 => b"01000_0000_01_000000000000", -- mul, gr0
 220 => b"00000_0000_00_000000001111", -- 15
 221 => b"00010_0000_00_000011110011", -- add, gr0, XPOS2
 222 => b"10000_0000_00_000000000000", -- tpoint, gr0
 223 => b"01111_0001_00_000000000000", -- tread, gr1
 224 => b"00011_0001_00_000011101100", -- sub, gr1, GRASS
 225 => b"00111_0000_01_000000000000", -- bne
 226 => b"00000_0000_00_000000000100", -- CONTROL_R
 227 => b"00010_1111_01_000000000000", -- add, gr15
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00100_0000_01_000000000000", -- jump
 230 => b"00000_0000_00_000000000100", -- CONTROL_R
 231 => b"00100_0000_01_000000000000", -- jump
 232 => b"00000_0000_00_000001001101", -- COUNT_R
 233 => b"00000_0000_00_000000000000", -- 0
 234 => b"00000_0000_00_000000000000", -- 0
 235 => b"00000_0000_00_000000000011", -- 3
 236 => b"00000_0000_00_000000000000", -- 0
 237 => b"00000_0000_00_000000000001", -- 1
 238 => b"00000_0000_00_000000000010", -- 2
 239 => b"00000_0000_00_000000000011", -- 3
 240 => b"00000_0000_00_000000000100", -- 4
 241 => b"00000_0000_00_000000000000", -- 0
 242 => b"00000_0000_00_000000000000", -- 0
 243 => b"00000_0000_00_000000000000", -- 0
 244 => b"00000_0000_00_000000000000", -- 0
 245 => b"00000_0000_00_000000000000", -- 0
 246 => b"00000_0000_00_000000000000", -- 0
 247 => b"00000_0000_00_000000000000", -- 0



   



    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


