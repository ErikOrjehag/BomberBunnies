library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr




    


    
0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000100010101", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011001011", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000001100110", -- TICKBOMBS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000001100", -- TICKEXPLOSIONS
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000000010", -- MAIN
  12 => b"00000_0000_00_000110110111", -- load, gr0, P1EXPLOSIONACTIVE
  13 => b"00011_0000_01_000000000000", -- sub, gr0
  14 => b"00000_0000_00_000000000001", -- 1
  15 => b"00111_0000_01_000000000000", -- bne
  16 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  17 => b"00000_0000_00_000110110110", -- load, gr0, P1EXPLOSIONTIME
  18 => b"00011_0000_01_000000000000", -- sub, gr0
  19 => b"00000_0000_00_000000000001", -- 1
  20 => b"00001_0000_10_000110110110", -- store, gr0, P1EXPLOSIONTIME
  21 => b"00000_0000_00_000110110110", -- load, gr0, P1EXPLOSIONTIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000000", -- 0
  24 => b"00111_0000_01_000000000000", -- bne
  25 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  26 => b"00000_0000_01_000000000000", -- load, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00001_0000_10_000110110111", -- store, gr0, P1EXPLOSIONACTIVE
  29 => b"00000_0010_00_000110111000", -- load, gr2, P1EXPLOSIONPOS
  30 => b"00000_0011_00_000111001001", -- load, gr3, GRASS
  31 => b"10000_0010_00_000000000000", -- tpoint, gr2
  32 => b"01110_0011_00_000000000000", -- twrite, gr3
  33 => b"00010_0010_01_000000000000", -- add, gr2
  34 => b"00000_0000_00_000000000001", -- 1
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01111_0000_00_000000000000", -- tread, gr0
  37 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  38 => b"00111_0000_01_000000000000", -- bne
  39 => b"00000_0000_00_000000110001", -- E1LEFT
  40 => b"01110_0011_00_000000000000", -- twrite, gr3
  41 => b"00010_0010_01_000000000000", -- add, gr2
  42 => b"00000_0000_00_000000000001", -- 1
  43 => b"10000_0010_00_000000000000", -- tpoint, gr2
  44 => b"01111_0000_00_000000000000", -- tread, gr0
  45 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  46 => b"00111_0000_01_000000000000", -- bne
  47 => b"00000_0000_00_000000110001", -- E1LEFT
  48 => b"01110_0011_00_000000000000", -- twrite, gr3
  49 => b"00000_0010_00_000110111000", -- load, gr2, P1EXPLOSIONPOS
  50 => b"00011_0010_01_000000000000", -- sub, gr2
  51 => b"00000_0000_00_000000000001", -- 1
  52 => b"10000_0010_00_000000000000", -- tpoint, gr2
  53 => b"01111_0000_00_000000000000", -- tread, gr0
  54 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  55 => b"00111_0000_01_000000000000", -- bne
  56 => b"00000_0000_00_000001000010", -- E1DOWN
  57 => b"01110_0011_00_000000000000", -- twrite, gr3
  58 => b"00011_0010_01_000000000000", -- sub, gr2
  59 => b"00000_0000_00_000000000001", -- 1
  60 => b"10000_0010_00_000000000000", -- tpoint, gr2
  61 => b"01111_0000_00_000000000000", -- tread, gr0
  62 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  63 => b"00111_0000_01_000000000000", -- bne
  64 => b"00000_0000_00_000001000010", -- E1DOWN
  65 => b"01110_0011_00_000000000000", -- twrite, gr3
  66 => b"00000_0010_00_000110111000", -- load, gr2, P1EXPLOSIONPOS
  67 => b"00010_0010_01_000000000000", -- add, gr2
  68 => b"00000_0000_00_000000001111", -- 15
  69 => b"10000_0010_00_000000000000", -- tpoint, gr2
  70 => b"01111_0000_00_000000000000", -- tread, gr0
  71 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  72 => b"00111_0000_01_000000000000", -- bne
  73 => b"00000_0000_00_000001010011", -- E1UP
  74 => b"01110_0011_00_000000000000", -- twrite, gr3
  75 => b"00010_0010_01_000000000000", -- add, gr2
  76 => b"00000_0000_00_000000001111", -- 15
  77 => b"10000_0010_00_000000000000", -- tpoint, gr2
  78 => b"01111_0000_00_000000000000", -- tread, gr0
  79 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  80 => b"00111_0000_01_000000000000", -- bne
  81 => b"00000_0000_00_000001010011", -- E1UP
  82 => b"01110_0011_00_000000000000", -- twrite, gr3
  83 => b"00000_0010_00_000110111000", -- load, gr2, P1EXPLOSIONPOS
  84 => b"00011_0010_01_000000000000", -- sub, gr2
  85 => b"00000_0000_00_000000001111", -- 15
  86 => b"10000_0010_00_000000000000", -- tpoint, gr2
  87 => b"01111_0000_00_000000000000", -- tread, gr0
  88 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  89 => b"00111_0000_01_000000000000", -- bne
  90 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  91 => b"01110_0011_00_000000000000", -- twrite, gr3
  92 => b"00011_0010_01_000000000000", -- sub, gr2
  93 => b"00000_0000_00_000000001111", -- 15
  94 => b"10000_0010_00_000000000000", -- tpoint, gr2
  95 => b"01111_0000_00_000000000000", -- tread, gr0
  96 => b"00011_0000_00_000111001100", -- sub, gr0, EXPLOSION
  97 => b"00111_0000_01_000000000000", -- bne
  98 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  99 => b"01110_0011_00_000000000000", -- twrite, gr3
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS_R
 102 => b"00000_0000_00_000110110101", -- load, gr0, P1BOMBACTIVE
 103 => b"00011_0000_01_000000000000", -- sub, gr0
 104 => b"00000_0000_00_000000000001", -- 1
 105 => b"00111_0000_01_000000000000", -- bne
 106 => b"00000_0000_00_000011001001", -- TICK2
 107 => b"00000_0000_00_000110110100", -- load, gr0, P1BOMBTIME
 108 => b"00011_0000_01_000000000000", -- sub, gr0
 109 => b"00000_0000_00_000000000001", -- 1
 110 => b"00001_0000_10_000110110100", -- store, gr0, P1BOMBTIME
 111 => b"00000_0000_01_000000000000", -- load, gr0
 112 => b"00000_0000_00_000000000000", -- 0
 113 => b"00011_0000_00_000110110100", -- sub, gr0, P1BOMBTIME
 114 => b"00110_0000_01_000000000000", -- beq
 115 => b"00000_0000_00_000001110110", -- EXPLODE1
 116 => b"00100_0000_01_000000000000", -- jump
 117 => b"00000_0000_00_000011001001", -- TICK2
 118 => b"00000_0000_00_000110110011", -- load, gr0, P1BOMBPOS
 119 => b"00001_0000_10_000110111000", -- store, gr0, P1EXPLOSIONPOS
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000001", -- 1
 122 => b"00001_0000_10_000110110111", -- store, gr0, P1EXPLOSIONACTIVE
 123 => b"00000_0000_01_000000000000", -- load, gr0
 124 => b"00000_0000_00_000000000010", -- 2
 125 => b"00001_0000_10_000110110110", -- store, gr0, P1EXPLOSIONTIME
 126 => b"00000_0000_00_000110111111", -- load, gr0, BOMBS1
 127 => b"00011_0000_01_000000000000", -- sub, gr0
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"00001_0000_10_000110111111", -- store, gr0, BOMBS1
 130 => b"00000_0010_00_000110110011", -- load, gr2, P1BOMBPOS
 131 => b"00000_0011_00_000111001100", -- load, gr3, EXPLOSION
 132 => b"10000_0010_00_000000000000", -- tpoint, gr2
 133 => b"01110_0011_00_000000000000", -- twrite, gr3
 134 => b"00010_0010_01_000000000000", -- add, gr2
 135 => b"00000_0000_00_000000000001", -- 1
 136 => b"10000_0010_00_000000000000", -- tpoint, gr2
 137 => b"01111_0000_00_000000000000", -- tread, gr0
 138 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 139 => b"00110_0000_01_000000000000", -- beq
 140 => b"00000_0000_00_000010010110", -- P1LEFT
 141 => b"01110_0011_00_000000000000", -- twrite, gr3
 142 => b"00010_0010_01_000000000000", -- add, gr2
 143 => b"00000_0000_00_000000000001", -- 1
 144 => b"10000_0010_00_000000000000", -- tpoint, gr2
 145 => b"01111_0000_00_000000000000", -- tread, gr0
 146 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 147 => b"00110_0000_01_000000000000", -- beq
 148 => b"00000_0000_00_000010010110", -- P1LEFT
 149 => b"01110_0011_00_000000000000", -- twrite, gr3
 150 => b"00000_0010_00_000110110011", -- load, gr2, P1BOMBPOS
 151 => b"00011_0010_01_000000000000", -- sub, gr2
 152 => b"00000_0000_00_000000000001", -- 1
 153 => b"10000_0010_00_000000000000", -- tpoint, gr2
 154 => b"01111_0000_00_000000000000", -- tread, gr0
 155 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 156 => b"00110_0000_01_000000000000", -- beq
 157 => b"00000_0000_00_000010100111", -- P1DOWN
 158 => b"01110_0011_00_000000000000", -- twrite, gr3
 159 => b"00011_0010_01_000000000000", -- sub, gr2
 160 => b"00000_0000_00_000000000001", -- 1
 161 => b"10000_0010_00_000000000000", -- tpoint, gr2
 162 => b"01111_0000_00_000000000000", -- tread, gr0
 163 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 164 => b"00110_0000_01_000000000000", -- beq
 165 => b"00000_0000_00_000010100111", -- P1DOWN
 166 => b"01110_0011_00_000000000000", -- twrite, gr3
 167 => b"00000_0010_00_000110110011", -- load, gr2, P1BOMBPOS
 168 => b"00010_0010_01_000000000000", -- add, gr2
 169 => b"00000_0000_00_000000001111", -- 15
 170 => b"10000_0010_00_000000000000", -- tpoint, gr2
 171 => b"01111_0000_00_000000000000", -- tread, gr0
 172 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 173 => b"00110_0000_01_000000000000", -- beq
 174 => b"00000_0000_00_000010111000", -- P1UP
 175 => b"01110_0011_00_000000000000", -- twrite, gr3
 176 => b"00010_0010_01_000000000000", -- add, gr2
 177 => b"00000_0000_00_000000001111", -- 15
 178 => b"10000_0010_00_000000000000", -- tpoint, gr2
 179 => b"01111_0000_00_000000000000", -- tread, gr0
 180 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 181 => b"00110_0000_01_000000000000", -- beq
 182 => b"00000_0000_00_000010111000", -- P1UP
 183 => b"01110_0011_00_000000000000", -- twrite, gr3
 184 => b"00000_0010_00_000110110011", -- load, gr2, P1BOMBPOS
 185 => b"00011_0010_01_000000000000", -- sub, gr2
 186 => b"00000_0000_00_000000001111", -- 15
 187 => b"10000_0010_00_000000000000", -- tpoint, gr2
 188 => b"01111_0000_00_000000000000", -- tread, gr0
 189 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 190 => b"00110_0000_01_000000000000", -- beq
 191 => b"00000_0000_00_000011001001", -- TICK2
 192 => b"01110_0011_00_000000000000", -- twrite, gr3
 193 => b"00011_0010_01_000000000000", -- sub, gr2
 194 => b"00000_0000_00_000000001111", -- 15
 195 => b"10000_0010_00_000000000000", -- tpoint, gr2
 196 => b"01111_0000_00_000000000000", -- tread, gr0
 197 => b"00011_0000_00_000111001010", -- sub, gr0, WALL
 198 => b"00110_0000_01_000000000000", -- beq
 199 => b"00000_0000_00_000011001001", -- TICK2
 200 => b"01110_0011_00_000000000000", -- twrite, gr3
 201 => b"00100_0000_01_000000000000", -- jump
 202 => b"00000_0000_00_000000001000", -- TICKBOMBS_R
 203 => b"10101_0000_01_000000000000", -- btn1
 204 => b"00000_0000_00_000011010001", -- BTN1
 205 => b"11010_0000_01_000000000000", -- btn2
 206 => b"00000_0000_00_000011110110", -- BTN2
 207 => b"00100_0000_01_000000000000", -- jump
 208 => b"00000_0000_00_000000000110", -- BUTTON_R
 209 => b"00000_0000_00_000110111111", -- load, gr0, BOMBS1
 210 => b"00011_0000_00_000111000001", -- sub, gr0, MAXBOMBS
 211 => b"00110_0000_01_000000000000", -- beq
 212 => b"00000_0000_00_000011001101", -- BTN1_R
 213 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 214 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 215 => b"00000_0000_00_000111000011", -- load, gr0, YPOS1
 216 => b"01000_0000_01_000000000000", -- mul, gr0
 217 => b"00000_0000_00_000000001111", -- 15
 218 => b"00010_0000_00_000111000010", -- add, gr0, XPOS1
 219 => b"10000_0000_00_000000000000", -- tpoint, gr0
 220 => b"01111_0001_00_000000000000", -- tread, gr1
 221 => b"00011_0001_00_000111001101", -- sub, gr1, EGG
 222 => b"00110_0000_01_000000000000", -- beq
 223 => b"00000_0000_00_000011001111", -- BTN2_R
 224 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 225 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 226 => b"00000_0011_00_000111000011", -- load, gr3, YPOS1
 227 => b"00000_0010_00_000111001101", -- load, gr2, EGG
 228 => b"01000_0011_01_000000000000", -- mul, gr3
 229 => b"00000_0000_00_000000001111", -- 15
 230 => b"00010_0011_00_000111000010", -- add, gr3, XPOS1
 231 => b"10000_0011_00_000000000000", -- tpoint, gr3
 232 => b"01110_0010_00_000000000000", -- twrite, gr2
 233 => b"00000_0000_01_000000000000", -- load, gr0
 234 => b"00000_0000_00_000000000001", -- 1
 235 => b"00001_0000_10_000110110101", -- store, gr0, P1BOMBACTIVE
 236 => b"00001_0011_10_000110110011", -- store, gr3, P1BOMBPOS
 237 => b"00000_0000_01_000000000000", -- load, gr0
 238 => b"00000_0000_00_000000010000", -- 16
 239 => b"00001_0000_10_000110110100", -- store, gr0, P1BOMBTIME
 240 => b"00000_0000_00_000110111111", -- load, gr0, BOMBS1
 241 => b"00010_0000_01_000000000000", -- add, gr0
 242 => b"00000_0000_00_000000000001", -- 1
 243 => b"00001_0000_10_000110111111", -- store, gr0, BOMBS1
 244 => b"00100_0000_01_000000000000", -- jump
 245 => b"00000_0000_00_000011001101", -- BTN1_R
 246 => b"00000_0000_00_000111000000", -- load, gr0, BOMBS2
 247 => b"00011_0000_00_000111000001", -- sub, gr0, MAXBOMBS
 248 => b"00110_0000_01_000000000000", -- beq
 249 => b"00000_0000_00_000011001111", -- BTN2_R
 250 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 251 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 252 => b"00000_0000_00_000111000101", -- load, gr0, YPOS2
 253 => b"01000_0000_01_000000000000", -- mul, gr0
 254 => b"00000_0000_00_000000001111", -- 15
 255 => b"00010_0000_00_000111000100", -- add, gr0, XPOS2
 256 => b"10000_0000_00_000000000000", -- tpoint, gr0
 257 => b"01111_0001_00_000000000000", -- tread, gr1
 258 => b"00011_0001_00_000111001101", -- sub, gr1, EGG
 259 => b"00110_0000_01_000000000000", -- beq
 260 => b"00000_0000_00_000011001111", -- BTN2_R
 261 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 262 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 263 => b"00000_0011_00_000111000101", -- load, gr3, YPOS2
 264 => b"00000_0010_00_000111001101", -- load, gr2, EGG
 265 => b"01000_0011_01_000000000000", -- mul, gr3
 266 => b"00000_0000_00_000000001111", -- 15
 267 => b"00010_0011_00_000111000100", -- add, gr3, XPOS2
 268 => b"10000_0011_00_000000000000", -- tpoint, gr3
 269 => b"01110_0010_00_000000000000", -- twrite, gr2
 270 => b"00000_0000_00_000111000000", -- load, gr0, BOMBS2
 271 => b"00010_0000_01_000000000000", -- add, gr0
 272 => b"00000_0000_00_000000000001", -- 1
 273 => b"00001_0000_10_000111000000", -- store, gr0, BOMBS2
 274 => b"00100_0000_01_000000000000", -- jump
 275 => b"00000_0000_00_000011001111", -- BTN2_R
 276 => b"00000_0000_00_000000000000", -- 0
 277 => b"00100_0000_01_000000000000", -- jump
 278 => b"00000_0000_00_000110110001", -- COUNT1
 279 => b"10001_0000_01_000000000000", -- joy1r
 280 => b"00000_0000_00_000100101001", -- P1R
 281 => b"10011_0000_01_000000000000", -- joy1l
 282 => b"00000_0000_00_000101001011", -- P1L
 283 => b"10010_0000_01_000000000000", -- joy1u
 284 => b"00000_0000_00_000100111010", -- P1U
 285 => b"10100_0000_01_000000000000", -- joy1d
 286 => b"00000_0000_00_000101011100", -- P1D
 287 => b"10110_0000_01_000000000000", -- joy2r
 288 => b"00000_0000_00_000101101101", -- P2R
 289 => b"11000_0000_01_000000000000", -- joy2l
 290 => b"00000_0000_00_000110001111", -- P2L
 291 => b"10111_0000_01_000000000000", -- joy2u
 292 => b"00000_0000_00_000101111110", -- P2U
 293 => b"11001_0000_01_000000000000", -- joy2d
 294 => b"00000_0000_00_000110100000", -- P2D
 295 => b"00100_0000_01_000000000000", -- jump
 296 => b"00000_0000_00_000000000100", -- CONTROL_R
 297 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 298 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 299 => b"00000_0000_00_000111000011", -- load, gr0, YPOS1
 300 => b"01000_0000_01_000000000000", -- mul, gr0
 301 => b"00000_0000_00_000000001111", -- 15
 302 => b"00010_0000_00_000111000010", -- add, gr0, XPOS1
 303 => b"00010_0000_01_000000000000", -- add, gr0
 304 => b"00000_0000_00_000000000001", -- 1
 305 => b"10000_0000_00_000000000000", -- tpoint, gr0
 306 => b"01111_0001_00_000000000000", -- tread, gr1
 307 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 308 => b"00111_0000_01_000000000000", -- bne
 309 => b"00000_0000_00_000100011011", -- J1
 310 => b"00010_1100_01_000000000000", -- add, gr12
 311 => b"00000_0000_00_000000000001", -- 1
 312 => b"00100_0000_01_000000000000", -- jump
 313 => b"00000_0000_00_000100011011", -- J1
 314 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 315 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 316 => b"00000_0000_00_000111000011", -- load, gr0, YPOS1
 317 => b"00011_0000_01_000000000000", -- sub, gr0
 318 => b"00000_0000_00_000000000001", -- 1
 319 => b"01000_0000_01_000000000000", -- mul, gr0
 320 => b"00000_0000_00_000000001111", -- 15
 321 => b"00010_0000_00_000111000010", -- add, gr0, XPOS1
 322 => b"10000_0000_00_000000000000", -- tpoint, gr0
 323 => b"01111_0001_00_000000000000", -- tread, gr1
 324 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 325 => b"00111_0000_01_000000000000", -- bne
 326 => b"00000_0000_00_000100011111", -- J2
 327 => b"00011_1101_01_000000000000", -- sub, gr13
 328 => b"00000_0000_00_000000000001", -- 1
 329 => b"00100_0000_01_000000000000", -- jump
 330 => b"00000_0000_00_000100011111", -- J2
 331 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 332 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 333 => b"00000_0000_00_000111000011", -- load, gr0, YPOS1
 334 => b"01000_0000_01_000000000000", -- mul, gr0
 335 => b"00000_0000_00_000000001111", -- 15
 336 => b"00010_0000_00_000111000010", -- add, gr0, XPOS1
 337 => b"00011_0000_01_000000000000", -- sub, gr0
 338 => b"00000_0000_00_000000000001", -- 1
 339 => b"10000_0000_00_000000000000", -- tpoint, gr0
 340 => b"01111_0001_00_000000000000", -- tread, gr1
 341 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 342 => b"00111_0000_01_000000000000", -- bne
 343 => b"00000_0000_00_000100011011", -- J1
 344 => b"00011_1100_01_000000000000", -- sub, gr12
 345 => b"00000_0000_00_000000000001", -- 1
 346 => b"00100_0000_01_000000000000", -- jump
 347 => b"00000_0000_00_000100011011", -- J1
 348 => b"00001_1100_10_000111000010", -- store, gr12, XPOS1
 349 => b"00001_1101_10_000111000011", -- store, gr13, YPOS1
 350 => b"00000_0000_00_000111000011", -- load, gr0, YPOS1
 351 => b"00010_0000_01_000000000000", -- add, gr0
 352 => b"00000_0000_00_000000000001", -- 1
 353 => b"01000_0000_01_000000000000", -- mul, gr0
 354 => b"00000_0000_00_000000001111", -- 15
 355 => b"00010_0000_00_000111000010", -- add, gr0, XPOS1
 356 => b"10000_0000_00_000000000000", -- tpoint, gr0
 357 => b"01111_0001_00_000000000000", -- tread, gr1
 358 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 359 => b"00111_0000_01_000000000000", -- bne
 360 => b"00000_0000_00_000100011111", -- J2
 361 => b"00010_1101_01_000000000000", -- add, gr13
 362 => b"00000_0000_00_000000000001", -- 1
 363 => b"00100_0000_01_000000000000", -- jump
 364 => b"00000_0000_00_000100011111", -- J2
 365 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 366 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 367 => b"00000_0000_00_000111000101", -- load, gr0, YPOS2
 368 => b"01000_0000_01_000000000000", -- mul, gr0
 369 => b"00000_0000_00_000000001111", -- 15
 370 => b"00010_0000_00_000111000100", -- add, gr0, XPOS2
 371 => b"00010_0000_01_000000000000", -- add, gr0
 372 => b"00000_0000_00_000000000001", -- 1
 373 => b"10000_0000_00_000000000000", -- tpoint, gr0
 374 => b"01111_0001_00_000000000000", -- tread, gr1
 375 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 376 => b"00111_0000_01_000000000000", -- bne
 377 => b"00000_0000_00_000100100011", -- J3
 378 => b"00010_1110_01_000000000000", -- add, gr14
 379 => b"00000_0000_00_000000000001", -- 1
 380 => b"00100_0000_01_000000000000", -- jump
 381 => b"00000_0000_00_000100100011", -- J3
 382 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 383 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 384 => b"00000_0000_00_000111000101", -- load, gr0, YPOS2
 385 => b"00011_0000_01_000000000000", -- sub, gr0
 386 => b"00000_0000_00_000000000001", -- 1
 387 => b"01000_0000_01_000000000000", -- mul, gr0
 388 => b"00000_0000_00_000000001111", -- 15
 389 => b"00010_0000_00_000111000100", -- add, gr0, XPOS2
 390 => b"10000_0000_00_000000000000", -- tpoint, gr0
 391 => b"01111_0001_00_000000000000", -- tread, gr1
 392 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 393 => b"00111_0000_01_000000000000", -- bne
 394 => b"00000_0000_00_000000000100", -- CONTROL_R
 395 => b"00011_1111_01_000000000000", -- sub, gr15
 396 => b"00000_0000_00_000000000001", -- 1
 397 => b"00100_0000_01_000000000000", -- jump
 398 => b"00000_0000_00_000000000100", -- CONTROL_R
 399 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 400 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 401 => b"00000_0000_00_000111000101", -- load, gr0, YPOS2
 402 => b"01000_0000_01_000000000000", -- mul, gr0
 403 => b"00000_0000_00_000000001111", -- 15
 404 => b"00010_0000_00_000111000100", -- add, gr0, XPOS2
 405 => b"00011_0000_01_000000000000", -- sub, gr0
 406 => b"00000_0000_00_000000000001", -- 1
 407 => b"10000_0000_00_000000000000", -- tpoint, gr0
 408 => b"01111_0001_00_000000000000", -- tread, gr1
 409 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 410 => b"00111_0000_01_000000000000", -- bne
 411 => b"00000_0000_00_000100100011", -- J3
 412 => b"00011_1110_01_000000000000", -- sub, gr14
 413 => b"00000_0000_00_000000000001", -- 1
 414 => b"00100_0000_01_000000000000", -- jump
 415 => b"00000_0000_00_000100100011", -- J3
 416 => b"00001_1110_10_000111000100", -- store, gr14, XPOS2
 417 => b"00001_1111_10_000111000101", -- store, gr15, YPOS2
 418 => b"00000_0000_00_000111000101", -- load, gr0, YPOS2
 419 => b"00010_0000_01_000000000000", -- add, gr0
 420 => b"00000_0000_00_000000000001", -- 1
 421 => b"01000_0000_01_000000000000", -- mul, gr0
 422 => b"00000_0000_00_000000001111", -- 15
 423 => b"00010_0000_00_000111000100", -- add, gr0, XPOS2
 424 => b"10000_0000_00_000000000000", -- tpoint, gr0
 425 => b"01111_0001_00_000000000000", -- tread, gr1
 426 => b"00011_0001_00_000111001001", -- sub, gr1, GRASS
 427 => b"00111_0000_01_000000000000", -- bne
 428 => b"00000_0000_00_000000000100", -- CONTROL_R
 429 => b"00010_1111_01_000000000000", -- add, gr15
 430 => b"00000_0000_00_000000000001", -- 1
 431 => b"00100_0000_01_000000000000", -- jump
 432 => b"00000_0000_00_000000000100", -- CONTROL_R
 433 => b"00100_0000_01_000000000000", -- jump
 434 => b"00000_0000_00_000100010111", -- COUNT_R
 435 => b"00000_0000_00_000000000000", -- 0
 436 => b"00000_0000_00_000000000000", -- 0
 437 => b"00000_0000_00_000000000000", -- 0
 438 => b"00000_0000_00_000000000000", -- 0
 439 => b"00000_0000_00_000000000000", -- 0
 440 => b"00000_0000_00_000000000000", -- 0
 441 => b"00000_0000_00_000000000000", -- 0
 442 => b"00000_0000_00_000000000000", -- 0
 443 => b"00000_0000_00_000000000000", -- 0
 444 => b"00000_0000_00_000000000000", -- 0
 445 => b"00000_0000_00_000000000000", -- 0
 446 => b"00000_0000_00_000000000000", -- 0
 447 => b"00000_0000_00_000000000000", -- 0
 448 => b"00000_0000_00_000000000000", -- 0
 449 => b"00000_0000_00_000000000001", -- 1
 450 => b"00000_0000_00_000000000000", -- 0
 451 => b"00000_0000_00_000000000000", -- 0
 452 => b"00000_0000_00_000000000000", -- 0
 453 => b"00000_0000_00_000000000000", -- 0
 454 => b"00000_0000_00_000000000000", -- 0
 455 => b"00000_0000_00_000000000000", -- 0
 456 => b"00000_0000_00_000000000000", -- 0
 457 => b"00000_0000_00_000000000000", -- 0
 458 => b"00000_0000_00_000000000001", -- 1
 459 => b"00000_0000_00_000000000010", -- 2
 460 => b"00000_0000_00_000000000011", -- 3
 461 => b"00000_0000_00_000000000100", -- 4



    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


