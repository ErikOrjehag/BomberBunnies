library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000111100111", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000110010110", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000011000110", -- TICKBOMBS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000001100", -- TICKEXPLOSIONS
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000000010", -- MAIN
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000000010010", -- BOOM1
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000001101100", -- BOOM2
  16 => b"00100_0000_01_000000000000", -- jump
  17 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS_R
  18 => b"00000_0000_00_001010001001", -- load, gr0, P1EXPLOSIONACTIVE
  19 => b"00011_0000_01_000000000000", -- sub, gr0
  20 => b"00000_0000_00_000000000001", -- 1
  21 => b"00111_0000_01_000000000000", -- bne
  22 => b"00000_0000_00_000000001110", -- BOOM1_R
  23 => b"00000_0000_00_001010001000", -- load, gr0, P1EXPLOSIONTIME
  24 => b"00011_0000_01_000000000000", -- sub, gr0
  25 => b"00000_0000_00_000000000001", -- 1
  26 => b"00001_0000_10_001010001000", -- store, gr0, P1EXPLOSIONTIME
  27 => b"00000_0000_00_001010001000", -- load, gr0, P1EXPLOSIONTIME
  28 => b"00011_0000_01_000000000000", -- sub, gr0
  29 => b"00000_0000_00_000000000000", -- 0
  30 => b"00111_0000_01_000000000000", -- bne
  31 => b"00000_0000_00_000000001110", -- BOOM1_R
  32 => b"00000_0000_01_000000000000", -- load, gr0
  33 => b"00000_0000_00_000000000000", -- 0
  34 => b"00001_0000_10_001010001001", -- store, gr0, P1EXPLOSIONACTIVE
  35 => b"00000_0010_00_001010001010", -- load, gr2, P1EXPLOSIONPOS
  36 => b"00000_0011_00_001010011011", -- load, gr3, GRASS
  37 => b"10000_0010_00_000000000000", -- tpoint, gr2
  38 => b"01110_0011_00_000000000000", -- twrite, gr3
  39 => b"00010_0010_01_000000000000", -- add, gr2
  40 => b"00000_0000_00_000000000001", -- 1
  41 => b"10000_0010_00_000000000000", -- tpoint, gr2
  42 => b"01111_0000_00_000000000000", -- tread, gr0
  43 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  44 => b"00111_0000_01_000000000000", -- bne
  45 => b"00000_0000_00_000000110111", -- E1LEFT
  46 => b"01110_0011_00_000000000000", -- twrite, gr3
  47 => b"00010_0010_01_000000000000", -- add, gr2
  48 => b"00000_0000_00_000000000001", -- 1
  49 => b"10000_0010_00_000000000000", -- tpoint, gr2
  50 => b"01111_0000_00_000000000000", -- tread, gr0
  51 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  52 => b"00111_0000_01_000000000000", -- bne
  53 => b"00000_0000_00_000000110111", -- E1LEFT
  54 => b"01110_0011_00_000000000000", -- twrite, gr3
  55 => b"00000_0010_00_001010001010", -- load, gr2, P1EXPLOSIONPOS
  56 => b"00011_0010_01_000000000000", -- sub, gr2
  57 => b"00000_0000_00_000000000001", -- 1
  58 => b"10000_0010_00_000000000000", -- tpoint, gr2
  59 => b"01111_0000_00_000000000000", -- tread, gr0
  60 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  61 => b"00111_0000_01_000000000000", -- bne
  62 => b"00000_0000_00_000001001000", -- E1DOWN
  63 => b"01110_0011_00_000000000000", -- twrite, gr3
  64 => b"00011_0010_01_000000000000", -- sub, gr2
  65 => b"00000_0000_00_000000000001", -- 1
  66 => b"10000_0010_00_000000000000", -- tpoint, gr2
  67 => b"01111_0000_00_000000000000", -- tread, gr0
  68 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  69 => b"00111_0000_01_000000000000", -- bne
  70 => b"00000_0000_00_000001001000", -- E1DOWN
  71 => b"01110_0011_00_000000000000", -- twrite, gr3
  72 => b"00000_0010_00_001010001010", -- load, gr2, P1EXPLOSIONPOS
  73 => b"00010_0010_01_000000000000", -- add, gr2
  74 => b"00000_0000_00_000000001111", -- 15
  75 => b"10000_0010_00_000000000000", -- tpoint, gr2
  76 => b"01111_0000_00_000000000000", -- tread, gr0
  77 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  78 => b"00111_0000_01_000000000000", -- bne
  79 => b"00000_0000_00_000001011001", -- E1UP
  80 => b"01110_0011_00_000000000000", -- twrite, gr3
  81 => b"00010_0010_01_000000000000", -- add, gr2
  82 => b"00000_0000_00_000000001111", -- 15
  83 => b"10000_0010_00_000000000000", -- tpoint, gr2
  84 => b"01111_0000_00_000000000000", -- tread, gr0
  85 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  86 => b"00111_0000_01_000000000000", -- bne
  87 => b"00000_0000_00_000001011001", -- E1UP
  88 => b"01110_0011_00_000000000000", -- twrite, gr3
  89 => b"00000_0010_00_001010001010", -- load, gr2, P1EXPLOSIONPOS
  90 => b"00011_0010_01_000000000000", -- sub, gr2
  91 => b"00000_0000_00_000000001111", -- 15
  92 => b"10000_0010_00_000000000000", -- tpoint, gr2
  93 => b"01111_0000_00_000000000000", -- tread, gr0
  94 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
  95 => b"00111_0000_01_000000000000", -- bne
  96 => b"00000_0000_00_000000001110", -- BOOM1_R
  97 => b"01110_0011_00_000000000000", -- twrite, gr3
  98 => b"00011_0010_01_000000000000", -- sub, gr2
  99 => b"00000_0000_00_000000001111", -- 15
 100 => b"10000_0010_00_000000000000", -- tpoint, gr2
 101 => b"01111_0000_00_000000000000", -- tread, gr0
 102 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 103 => b"00111_0000_01_000000000000", -- bne
 104 => b"00000_0000_00_000000001110", -- BOOM1_R
 105 => b"01110_0011_00_000000000000", -- twrite, gr3
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000000001110", -- BOOM1_R
 108 => b"00000_0000_00_001010001111", -- load, gr0, P2EXPLOSIONACTIVE
 109 => b"00011_0000_01_000000000000", -- sub, gr0
 110 => b"00000_0000_00_000000000001", -- 1
 111 => b"00111_0000_01_000000000000", -- bne
 112 => b"00000_0000_00_000000010000", -- BOOM2_R
 113 => b"00000_0000_00_001010001110", -- load, gr0, P2EXPLOSIONTIME
 114 => b"00011_0000_01_000000000000", -- sub, gr0
 115 => b"00000_0000_00_000000000001", -- 1
 116 => b"00001_0000_10_001010001110", -- store, gr0, P2EXPLOSIONTIME
 117 => b"00000_0000_00_001010001110", -- load, gr0, P2EXPLOSIONTIME
 118 => b"00011_0000_01_000000000000", -- sub, gr0
 119 => b"00000_0000_00_000000000000", -- 0
 120 => b"00111_0000_01_000000000000", -- bne
 121 => b"00000_0000_00_000000010000", -- BOOM2_R
 122 => b"00000_0000_01_000000000000", -- load, gr0
 123 => b"00000_0000_00_000000000000", -- 0
 124 => b"00001_0000_10_001010001111", -- store, gr0, P2EXPLOSIONACTIVE
 125 => b"00000_0010_00_001010010000", -- load, gr2, P2EXPLOSIONPOS
 126 => b"00000_0011_00_001010011011", -- load, gr3, GRASS
 127 => b"10000_0010_00_000000000000", -- tpoint, gr2
 128 => b"01110_0011_00_000000000000", -- twrite, gr3
 129 => b"00010_0010_01_000000000000", -- add, gr2
 130 => b"00000_0000_00_000000000001", -- 1
 131 => b"10000_0010_00_000000000000", -- tpoint, gr2
 132 => b"01111_0000_00_000000000000", -- tread, gr0
 133 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 134 => b"00111_0000_01_000000000000", -- bne
 135 => b"00000_0000_00_000010010001", -- E2LEFT
 136 => b"01110_0011_00_000000000000", -- twrite, gr3
 137 => b"00010_0010_01_000000000000", -- add, gr2
 138 => b"00000_0000_00_000000000001", -- 1
 139 => b"10000_0010_00_000000000000", -- tpoint, gr2
 140 => b"01111_0000_00_000000000000", -- tread, gr0
 141 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 142 => b"00111_0000_01_000000000000", -- bne
 143 => b"00000_0000_00_000010010001", -- E2LEFT
 144 => b"01110_0011_00_000000000000", -- twrite, gr3
 145 => b"00000_0010_00_001010010000", -- load, gr2, P2EXPLOSIONPOS
 146 => b"00011_0010_01_000000000000", -- sub, gr2
 147 => b"00000_0000_00_000000000001", -- 1
 148 => b"10000_0010_00_000000000000", -- tpoint, gr2
 149 => b"01111_0000_00_000000000000", -- tread, gr0
 150 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 151 => b"00111_0000_01_000000000000", -- bne
 152 => b"00000_0000_00_000010100010", -- E2DOWN
 153 => b"01110_0011_00_000000000000", -- twrite, gr3
 154 => b"00011_0010_01_000000000000", -- sub, gr2
 155 => b"00000_0000_00_000000000001", -- 1
 156 => b"10000_0010_00_000000000000", -- tpoint, gr2
 157 => b"01111_0000_00_000000000000", -- tread, gr0
 158 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 159 => b"00111_0000_01_000000000000", -- bne
 160 => b"00000_0000_00_000010100010", -- E2DOWN
 161 => b"01110_0011_00_000000000000", -- twrite, gr3
 162 => b"00000_0010_00_001010010000", -- load, gr2, P2EXPLOSIONPOS
 163 => b"00010_0010_01_000000000000", -- add, gr2
 164 => b"00000_0000_00_000000001111", -- 15
 165 => b"10000_0010_00_000000000000", -- tpoint, gr2
 166 => b"01111_0000_00_000000000000", -- tread, gr0
 167 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 168 => b"00111_0000_01_000000000000", -- bne
 169 => b"00000_0000_00_000010110011", -- E2UP
 170 => b"01110_0011_00_000000000000", -- twrite, gr3
 171 => b"00010_0010_01_000000000000", -- add, gr2
 172 => b"00000_0000_00_000000001111", -- 15
 173 => b"10000_0010_00_000000000000", -- tpoint, gr2
 174 => b"01111_0000_00_000000000000", -- tread, gr0
 175 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 176 => b"00111_0000_01_000000000000", -- bne
 177 => b"00000_0000_00_000010110011", -- E2UP
 178 => b"01110_0011_00_000000000000", -- twrite, gr3
 179 => b"00000_0010_00_001010010000", -- load, gr2, P2EXPLOSIONPOS
 180 => b"00011_0010_01_000000000000", -- sub, gr2
 181 => b"00000_0000_00_000000001111", -- 15
 182 => b"10000_0010_00_000000000000", -- tpoint, gr2
 183 => b"01111_0000_00_000000000000", -- tread, gr0
 184 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 185 => b"00111_0000_01_000000000000", -- bne
 186 => b"00000_0000_00_000000010000", -- BOOM2_R
 187 => b"01110_0011_00_000000000000", -- twrite, gr3
 188 => b"00011_0010_01_000000000000", -- sub, gr2
 189 => b"00000_0000_00_000000001111", -- 15
 190 => b"10000_0010_00_000000000000", -- tpoint, gr2
 191 => b"01111_0000_00_000000000000", -- tread, gr0
 192 => b"00011_0000_00_001010011110", -- sub, gr0, EXPLOSION
 193 => b"00111_0000_01_000000000000", -- bne
 194 => b"00000_0000_00_000000010000", -- BOOM2_R
 195 => b"01110_0011_00_000000000000", -- twrite, gr3
 196 => b"00100_0000_01_000000000000", -- jump
 197 => b"00000_0000_00_000000010000", -- BOOM2_R
 198 => b"00100_0000_01_000000000000", -- jump
 199 => b"00000_0000_00_000011001100", -- TICKBOMB1
 200 => b"00100_0000_01_000000000000", -- jump
 201 => b"00000_0000_00_000100110001", -- TICKBOMB2
 202 => b"00100_0000_01_000000000000", -- jump
 203 => b"00000_0000_00_000000001000", -- TICKBOMBS_R
 204 => b"00000_0000_00_001010000111", -- load, gr0, P1BOMBACTIVE
 205 => b"00011_0000_01_000000000000", -- sub, gr0
 206 => b"00000_0000_00_000000000001", -- 1
 207 => b"00111_0000_01_000000000000", -- bne
 208 => b"00000_0000_00_000011001000", -- TICKBOMB1_R
 209 => b"00000_0000_00_001010000110", -- load, gr0, P1BOMBTIME
 210 => b"00011_0000_01_000000000000", -- sub, gr0
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00001_0000_10_001010000110", -- store, gr0, P1BOMBTIME
 213 => b"00000_0000_01_000000000000", -- load, gr0
 214 => b"00000_0000_00_000000000000", -- 0
 215 => b"00011_0000_00_001010000110", -- sub, gr0, P1BOMBTIME
 216 => b"00110_0000_01_000000000000", -- beq
 217 => b"00000_0000_00_000011011100", -- EXPLODE1
 218 => b"00100_0000_01_000000000000", -- jump
 219 => b"00000_0000_00_000011001000", -- TICKBOMB1_R
 220 => b"00000_0000_00_001010000101", -- load, gr0, P1BOMBPOS
 221 => b"00001_0000_10_001010001010", -- store, gr0, P1EXPLOSIONPOS
 222 => b"00000_0000_01_000000000000", -- load, gr0
 223 => b"00000_0000_00_000000000001", -- 1
 224 => b"00001_0000_10_001010001001", -- store, gr0, P1EXPLOSIONACTIVE
 225 => b"00000_0000_01_000000000000", -- load, gr0
 226 => b"00000_0000_00_000000000010", -- 2
 227 => b"00001_0000_10_001010001000", -- store, gr0, P1EXPLOSIONTIME
 228 => b"00000_0000_00_001010010001", -- load, gr0, BOMBS1
 229 => b"00011_0000_01_000000000000", -- sub, gr0
 230 => b"00000_0000_00_000000000001", -- 1
 231 => b"00001_0000_10_001010010001", -- store, gr0, BOMBS1
 232 => b"00000_0010_00_001010000101", -- load, gr2, P1BOMBPOS
 233 => b"00000_0011_00_001010011110", -- load, gr3, EXPLOSION
 234 => b"10000_0010_00_000000000000", -- tpoint, gr2
 235 => b"01110_0011_00_000000000000", -- twrite, gr3
 236 => b"00010_0010_01_000000000000", -- add, gr2
 237 => b"00000_0000_00_000000000001", -- 1
 238 => b"10000_0010_00_000000000000", -- tpoint, gr2
 239 => b"01111_0000_00_000000000000", -- tread, gr0
 240 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 241 => b"00110_0000_01_000000000000", -- beq
 242 => b"00000_0000_00_000011111100", -- P1LEFT
 243 => b"01110_0011_00_000000000000", -- twrite, gr3
 244 => b"00010_0010_01_000000000000", -- add, gr2
 245 => b"00000_0000_00_000000000001", -- 1
 246 => b"10000_0010_00_000000000000", -- tpoint, gr2
 247 => b"01111_0000_00_000000000000", -- tread, gr0
 248 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 249 => b"00110_0000_01_000000000000", -- beq
 250 => b"00000_0000_00_000011111100", -- P1LEFT
 251 => b"01110_0011_00_000000000000", -- twrite, gr3
 252 => b"00000_0010_00_001010000101", -- load, gr2, P1BOMBPOS
 253 => b"00011_0010_01_000000000000", -- sub, gr2
 254 => b"00000_0000_00_000000000001", -- 1
 255 => b"10000_0010_00_000000000000", -- tpoint, gr2
 256 => b"01111_0000_00_000000000000", -- tread, gr0
 257 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 258 => b"00110_0000_01_000000000000", -- beq
 259 => b"00000_0000_00_000100001101", -- P1DOWN
 260 => b"01110_0011_00_000000000000", -- twrite, gr3
 261 => b"00011_0010_01_000000000000", -- sub, gr2
 262 => b"00000_0000_00_000000000001", -- 1
 263 => b"10000_0010_00_000000000000", -- tpoint, gr2
 264 => b"01111_0000_00_000000000000", -- tread, gr0
 265 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 266 => b"00110_0000_01_000000000000", -- beq
 267 => b"00000_0000_00_000100001101", -- P1DOWN
 268 => b"01110_0011_00_000000000000", -- twrite, gr3
 269 => b"00000_0010_00_001010000101", -- load, gr2, P1BOMBPOS
 270 => b"00010_0010_01_000000000000", -- add, gr2
 271 => b"00000_0000_00_000000001111", -- 15
 272 => b"10000_0010_00_000000000000", -- tpoint, gr2
 273 => b"01111_0000_00_000000000000", -- tread, gr0
 274 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 275 => b"00110_0000_01_000000000000", -- beq
 276 => b"00000_0000_00_000100011110", -- P1UP
 277 => b"01110_0011_00_000000000000", -- twrite, gr3
 278 => b"00010_0010_01_000000000000", -- add, gr2
 279 => b"00000_0000_00_000000001111", -- 15
 280 => b"10000_0010_00_000000000000", -- tpoint, gr2
 281 => b"01111_0000_00_000000000000", -- tread, gr0
 282 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 283 => b"00110_0000_01_000000000000", -- beq
 284 => b"00000_0000_00_000100011110", -- P1UP
 285 => b"01110_0011_00_000000000000", -- twrite, gr3
 286 => b"00000_0010_00_001010000101", -- load, gr2, P1BOMBPOS
 287 => b"00011_0010_01_000000000000", -- sub, gr2
 288 => b"00000_0000_00_000000001111", -- 15
 289 => b"10000_0010_00_000000000000", -- tpoint, gr2
 290 => b"01111_0000_00_000000000000", -- tread, gr0
 291 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 292 => b"00110_0000_01_000000000000", -- beq
 293 => b"00000_0000_00_000011001000", -- TICKBOMB1_R
 294 => b"01110_0011_00_000000000000", -- twrite, gr3
 295 => b"00011_0010_01_000000000000", -- sub, gr2
 296 => b"00000_0000_00_000000001111", -- 15
 297 => b"10000_0010_00_000000000000", -- tpoint, gr2
 298 => b"01111_0000_00_000000000000", -- tread, gr0
 299 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 300 => b"00110_0000_01_000000000000", -- beq
 301 => b"00000_0000_00_000011001000", -- TICKBOMB1_R
 302 => b"01110_0011_00_000000000000", -- twrite, gr3
 303 => b"00100_0000_01_000000000000", -- jump
 304 => b"00000_0000_00_000011001000", -- TICKBOMB1_R
 305 => b"00000_0000_00_001010001101", -- load, gr0, P2BOMBACTIVE
 306 => b"00011_0000_01_000000000000", -- sub, gr0
 307 => b"00000_0000_00_000000000001", -- 1
 308 => b"00111_0000_01_000000000000", -- bne
 309 => b"00000_0000_00_000011001010", -- TICKBOMB2_R
 310 => b"00000_0000_00_001010001100", -- load, gr0, P2BOMBTIME
 311 => b"00011_0000_01_000000000000", -- sub, gr0
 312 => b"00000_0000_00_000000000001", -- 1
 313 => b"00001_0000_10_001010001100", -- store, gr0, P2BOMBTIME
 314 => b"00000_0000_01_000000000000", -- load, gr0
 315 => b"00000_0000_00_000000000000", -- 0
 316 => b"00011_0000_00_001010001100", -- sub, gr0, P2BOMBTIME
 317 => b"00110_0000_01_000000000000", -- beq
 318 => b"00000_0000_00_000101000001", -- EXPLODE2
 319 => b"00100_0000_01_000000000000", -- jump
 320 => b"00000_0000_00_000011001010", -- TICKBOMB2_R
 321 => b"00000_0000_00_001010001011", -- load, gr0, P2BOMBPOS
 322 => b"00001_0000_10_001010010000", -- store, gr0, P2EXPLOSIONPOS
 323 => b"00000_0000_01_000000000000", -- load, gr0
 324 => b"00000_0000_00_000000000001", -- 1
 325 => b"00001_0000_10_001010001111", -- store, gr0, P2EXPLOSIONACTIVE
 326 => b"00000_0000_01_000000000000", -- load, gr0
 327 => b"00000_0000_00_000000000010", -- 2
 328 => b"00001_0000_10_001010001110", -- store, gr0, P2EXPLOSIONTIME
 329 => b"00000_0000_00_001010010010", -- load, gr0, BOMBS2
 330 => b"00011_0000_01_000000000000", -- sub, gr0
 331 => b"00000_0000_00_000000000001", -- 1
 332 => b"00001_0000_10_001010010010", -- store, gr0, BOMBS2
 333 => b"00000_0010_00_001010001011", -- load, gr2, P2BOMBPOS
 334 => b"00000_0011_00_001010011110", -- load, gr3, EXPLOSION
 335 => b"10000_0010_00_000000000000", -- tpoint, gr2
 336 => b"01110_0011_00_000000000000", -- twrite, gr3
 337 => b"00010_0010_01_000000000000", -- add, gr2
 338 => b"00000_0000_00_000000000001", -- 1
 339 => b"10000_0010_00_000000000000", -- tpoint, gr2
 340 => b"01111_0000_00_000000000000", -- tread, gr0
 341 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 342 => b"00110_0000_01_000000000000", -- beq
 343 => b"00000_0000_00_000101100001", -- P2LEFT
 344 => b"01110_0011_00_000000000000", -- twrite, gr3
 345 => b"00010_0010_01_000000000000", -- add, gr2
 346 => b"00000_0000_00_000000000001", -- 1
 347 => b"10000_0010_00_000000000000", -- tpoint, gr2
 348 => b"01111_0000_00_000000000000", -- tread, gr0
 349 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 350 => b"00110_0000_01_000000000000", -- beq
 351 => b"00000_0000_00_000101100001", -- P2LEFT
 352 => b"01110_0011_00_000000000000", -- twrite, gr3
 353 => b"00000_0010_00_001010001011", -- load, gr2, P2BOMBPOS
 354 => b"00011_0010_01_000000000000", -- sub, gr2
 355 => b"00000_0000_00_000000000001", -- 1
 356 => b"10000_0010_00_000000000000", -- tpoint, gr2
 357 => b"01111_0000_00_000000000000", -- tread, gr0
 358 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 359 => b"00110_0000_01_000000000000", -- beq
 360 => b"00000_0000_00_000101110010", -- P2DOWN
 361 => b"01110_0011_00_000000000000", -- twrite, gr3
 362 => b"00011_0010_01_000000000000", -- sub, gr2
 363 => b"00000_0000_00_000000000001", -- 1
 364 => b"10000_0010_00_000000000000", -- tpoint, gr2
 365 => b"01111_0000_00_000000000000", -- tread, gr0
 366 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 367 => b"00110_0000_01_000000000000", -- beq
 368 => b"00000_0000_00_000101110010", -- P2DOWN
 369 => b"01110_0011_00_000000000000", -- twrite, gr3
 370 => b"00000_0010_00_001010001011", -- load, gr2, P2BOMBPOS
 371 => b"00010_0010_01_000000000000", -- add, gr2
 372 => b"00000_0000_00_000000001111", -- 15
 373 => b"10000_0010_00_000000000000", -- tpoint, gr2
 374 => b"01111_0000_00_000000000000", -- tread, gr0
 375 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 376 => b"00110_0000_01_000000000000", -- beq
 377 => b"00000_0000_00_000110000011", -- P2UP
 378 => b"01110_0011_00_000000000000", -- twrite, gr3
 379 => b"00010_0010_01_000000000000", -- add, gr2
 380 => b"00000_0000_00_000000001111", -- 15
 381 => b"10000_0010_00_000000000000", -- tpoint, gr2
 382 => b"01111_0000_00_000000000000", -- tread, gr0
 383 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 384 => b"00110_0000_01_000000000000", -- beq
 385 => b"00000_0000_00_000110000011", -- P2UP
 386 => b"01110_0011_00_000000000000", -- twrite, gr3
 387 => b"00000_0010_00_001010001011", -- load, gr2, P2BOMBPOS
 388 => b"00011_0010_01_000000000000", -- sub, gr2
 389 => b"00000_0000_00_000000001111", -- 15
 390 => b"10000_0010_00_000000000000", -- tpoint, gr2
 391 => b"01111_0000_00_000000000000", -- tread, gr0
 392 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 393 => b"00110_0000_01_000000000000", -- beq
 394 => b"00000_0000_00_000011001010", -- TICKBOMB2_R
 395 => b"01110_0011_00_000000000000", -- twrite, gr3
 396 => b"00011_0010_01_000000000000", -- sub, gr2
 397 => b"00000_0000_00_000000001111", -- 15
 398 => b"10000_0010_00_000000000000", -- tpoint, gr2
 399 => b"01111_0000_00_000000000000", -- tread, gr0
 400 => b"00011_0000_00_001010011100", -- sub, gr0, WALL
 401 => b"00110_0000_01_000000000000", -- beq
 402 => b"00000_0000_00_000011001010", -- TICKBOMB2_R
 403 => b"01110_0011_00_000000000000", -- twrite, gr3
 404 => b"00100_0000_01_000000000000", -- jump
 405 => b"00000_0000_00_000011001010", -- TICKBOMB2_R
 406 => b"10101_0000_01_000000000000", -- btn1
 407 => b"00000_0000_00_000110011100", -- BTN1
 408 => b"11010_0000_01_000000000000", -- btn2
 409 => b"00000_0000_00_000111000001", -- BTN2
 410 => b"00100_0000_01_000000000000", -- jump
 411 => b"00000_0000_00_000000000110", -- BUTTON_R
 412 => b"00000_0000_00_001010010001", -- load, gr0, BOMBS1
 413 => b"00011_0000_00_001010010011", -- sub, gr0, MAXBOMBS
 414 => b"00110_0000_01_000000000000", -- beq
 415 => b"00000_0000_00_000110011000", -- BTN1_R
 416 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 417 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 418 => b"00000_0000_00_001010010101", -- load, gr0, YPOS1
 419 => b"01000_0000_01_000000000000", -- mul, gr0
 420 => b"00000_0000_00_000000001111", -- 15
 421 => b"00010_0000_00_001010010100", -- add, gr0, XPOS1
 422 => b"10000_0000_00_000000000000", -- tpoint, gr0
 423 => b"01111_0001_00_000000000000", -- tread, gr1
 424 => b"00011_0001_00_001010011111", -- sub, gr1, EGG
 425 => b"00110_0000_01_000000000000", -- beq
 426 => b"00000_0000_00_000110011000", -- BTN1_R
 427 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 428 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 429 => b"00000_0011_00_001010010101", -- load, gr3, YPOS1
 430 => b"00000_0010_00_001010011111", -- load, gr2, EGG
 431 => b"01000_0011_01_000000000000", -- mul, gr3
 432 => b"00000_0000_00_000000001111", -- 15
 433 => b"00010_0011_00_001010010100", -- add, gr3, XPOS1
 434 => b"10000_0011_00_000000000000", -- tpoint, gr3
 435 => b"01110_0010_00_000000000000", -- twrite, gr2
 436 => b"00000_0000_01_000000000000", -- load, gr0
 437 => b"00000_0000_00_000000000001", -- 1
 438 => b"00001_0000_10_001010000111", -- store, gr0, P1BOMBACTIVE
 439 => b"00001_0011_10_001010000101", -- store, gr3, P1BOMBPOS
 440 => b"00000_0000_01_000000000000", -- load, gr0
 441 => b"00000_0000_00_000000010000", -- 16
 442 => b"00001_0000_10_001010000110", -- store, gr0, P1BOMBTIME
 443 => b"00000_0000_00_001010010001", -- load, gr0, BOMBS1
 444 => b"00010_0000_01_000000000000", -- add, gr0
 445 => b"00000_0000_00_000000000001", -- 1
 446 => b"00001_0000_10_001010010001", -- store, gr0, BOMBS1
 447 => b"00100_0000_01_000000000000", -- jump
 448 => b"00000_0000_00_000110011000", -- BTN1_R
 449 => b"00000_0000_00_001010010010", -- load, gr0, BOMBS2
 450 => b"00011_0000_00_001010010011", -- sub, gr0, MAXBOMBS
 451 => b"00110_0000_01_000000000000", -- beq
 452 => b"00000_0000_00_000110011010", -- BTN2_R
 453 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 454 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 455 => b"00000_0000_00_001010010111", -- load, gr0, YPOS2
 456 => b"01000_0000_01_000000000000", -- mul, gr0
 457 => b"00000_0000_00_000000001111", -- 15
 458 => b"00010_0000_00_001010010110", -- add, gr0, XPOS2
 459 => b"10000_0000_00_000000000000", -- tpoint, gr0
 460 => b"01111_0001_00_000000000000", -- tread, gr1
 461 => b"00011_0001_00_001010011111", -- sub, gr1, EGG
 462 => b"00110_0000_01_000000000000", -- beq
 463 => b"00000_0000_00_000110011010", -- BTN2_R
 464 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 465 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 466 => b"00000_0011_00_001010010111", -- load, gr3, YPOS2
 467 => b"00000_0010_00_001010011111", -- load, gr2, EGG
 468 => b"01000_0011_01_000000000000", -- mul, gr3
 469 => b"00000_0000_00_000000001111", -- 15
 470 => b"00010_0011_00_001010010110", -- add, gr3, XPOS2
 471 => b"10000_0011_00_000000000000", -- tpoint, gr3
 472 => b"01110_0010_00_000000000000", -- twrite, gr2
 473 => b"00000_0000_01_000000000000", -- load, gr0
 474 => b"00000_0000_00_000000000001", -- 1
 475 => b"00001_0000_10_001010001101", -- store, gr0, P2BOMBACTIVE
 476 => b"00001_0011_10_001010001011", -- store, gr3, P2BOMBPOS
 477 => b"00000_0000_01_000000000000", -- load, gr0
 478 => b"00000_0000_00_000000010000", -- 16
 479 => b"00001_0000_10_001010001100", -- store, gr0, P2BOMBTIME
 480 => b"00000_0000_00_001010010010", -- load, gr0, BOMBS2
 481 => b"00010_0000_01_000000000000", -- add, gr0
 482 => b"00000_0000_00_000000000001", -- 1
 483 => b"00001_0000_10_001010010010", -- store, gr0, BOMBS2
 484 => b"00100_0000_01_000000000000", -- jump
 485 => b"00000_0000_00_000110011010", -- BTN2_R
 486 => b"00000_0000_00_000000000000", -- 0
 487 => b"00100_0000_01_000000000000", -- jump
 488 => b"00000_0000_00_001010000011", -- COUNT1
 489 => b"10001_0000_01_000000000000", -- joy1r
 490 => b"00000_0000_00_000111111011", -- P1R
 491 => b"10011_0000_01_000000000000", -- joy1l
 492 => b"00000_0000_00_001000011101", -- P1L
 493 => b"10010_0000_01_000000000000", -- joy1u
 494 => b"00000_0000_00_001000001100", -- P1U
 495 => b"10100_0000_01_000000000000", -- joy1d
 496 => b"00000_0000_00_001000101110", -- P1D
 497 => b"10110_0000_01_000000000000", -- joy2r
 498 => b"00000_0000_00_001000111111", -- P2R
 499 => b"11000_0000_01_000000000000", -- joy2l
 500 => b"00000_0000_00_001001100001", -- P2L
 501 => b"10111_0000_01_000000000000", -- joy2u
 502 => b"00000_0000_00_001001010000", -- P2U
 503 => b"11001_0000_01_000000000000", -- joy2d
 504 => b"00000_0000_00_001001110010", -- P2D
 505 => b"00100_0000_01_000000000000", -- jump
 506 => b"00000_0000_00_000000000100", -- CONTROL_R
 507 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 508 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 509 => b"00000_0000_00_001010010101", -- load, gr0, YPOS1
 510 => b"01000_0000_01_000000000000", -- mul, gr0
 511 => b"00000_0000_00_000000001111", -- 15
 512 => b"00010_0000_00_001010010100", -- add, gr0, XPOS1
 513 => b"00010_0000_01_000000000000", -- add, gr0
 514 => b"00000_0000_00_000000000001", -- 1
 515 => b"10000_0000_00_000000000000", -- tpoint, gr0
 516 => b"01111_0001_00_000000000000", -- tread, gr1
 517 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 518 => b"00111_0000_01_000000000000", -- bne
 519 => b"00000_0000_00_000111101101", -- J1
 520 => b"00010_1100_01_000000000000", -- add, gr12
 521 => b"00000_0000_00_000000000001", -- 1
 522 => b"00100_0000_01_000000000000", -- jump
 523 => b"00000_0000_00_000111101101", -- J1
 524 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 525 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 526 => b"00000_0000_00_001010010101", -- load, gr0, YPOS1
 527 => b"00011_0000_01_000000000000", -- sub, gr0
 528 => b"00000_0000_00_000000000001", -- 1
 529 => b"01000_0000_01_000000000000", -- mul, gr0
 530 => b"00000_0000_00_000000001111", -- 15
 531 => b"00010_0000_00_001010010100", -- add, gr0, XPOS1
 532 => b"10000_0000_00_000000000000", -- tpoint, gr0
 533 => b"01111_0001_00_000000000000", -- tread, gr1
 534 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 535 => b"00111_0000_01_000000000000", -- bne
 536 => b"00000_0000_00_000111110001", -- J2
 537 => b"00011_1101_01_000000000000", -- sub, gr13
 538 => b"00000_0000_00_000000000001", -- 1
 539 => b"00100_0000_01_000000000000", -- jump
 540 => b"00000_0000_00_000111110001", -- J2
 541 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 542 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 543 => b"00000_0000_00_001010010101", -- load, gr0, YPOS1
 544 => b"01000_0000_01_000000000000", -- mul, gr0
 545 => b"00000_0000_00_000000001111", -- 15
 546 => b"00010_0000_00_001010010100", -- add, gr0, XPOS1
 547 => b"00011_0000_01_000000000000", -- sub, gr0
 548 => b"00000_0000_00_000000000001", -- 1
 549 => b"10000_0000_00_000000000000", -- tpoint, gr0
 550 => b"01111_0001_00_000000000000", -- tread, gr1
 551 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 552 => b"00111_0000_01_000000000000", -- bne
 553 => b"00000_0000_00_000111101101", -- J1
 554 => b"00011_1100_01_000000000000", -- sub, gr12
 555 => b"00000_0000_00_000000000001", -- 1
 556 => b"00100_0000_01_000000000000", -- jump
 557 => b"00000_0000_00_000111101101", -- J1
 558 => b"00001_1100_10_001010010100", -- store, gr12, XPOS1
 559 => b"00001_1101_10_001010010101", -- store, gr13, YPOS1
 560 => b"00000_0000_00_001010010101", -- load, gr0, YPOS1
 561 => b"00010_0000_01_000000000000", -- add, gr0
 562 => b"00000_0000_00_000000000001", -- 1
 563 => b"01000_0000_01_000000000000", -- mul, gr0
 564 => b"00000_0000_00_000000001111", -- 15
 565 => b"00010_0000_00_001010010100", -- add, gr0, XPOS1
 566 => b"10000_0000_00_000000000000", -- tpoint, gr0
 567 => b"01111_0001_00_000000000000", -- tread, gr1
 568 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 569 => b"00111_0000_01_000000000000", -- bne
 570 => b"00000_0000_00_000111110001", -- J2
 571 => b"00010_1101_01_000000000000", -- add, gr13
 572 => b"00000_0000_00_000000000001", -- 1
 573 => b"00100_0000_01_000000000000", -- jump
 574 => b"00000_0000_00_000111110001", -- J2
 575 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 576 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 577 => b"00000_0000_00_001010010111", -- load, gr0, YPOS2
 578 => b"01000_0000_01_000000000000", -- mul, gr0
 579 => b"00000_0000_00_000000001111", -- 15
 580 => b"00010_0000_00_001010010110", -- add, gr0, XPOS2
 581 => b"00010_0000_01_000000000000", -- add, gr0
 582 => b"00000_0000_00_000000000001", -- 1
 583 => b"10000_0000_00_000000000000", -- tpoint, gr0
 584 => b"01111_0001_00_000000000000", -- tread, gr1
 585 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 586 => b"00111_0000_01_000000000000", -- bne
 587 => b"00000_0000_00_000111110101", -- J3
 588 => b"00010_1110_01_000000000000", -- add, gr14
 589 => b"00000_0000_00_000000000001", -- 1
 590 => b"00100_0000_01_000000000000", -- jump
 591 => b"00000_0000_00_000111110101", -- J3
 592 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 593 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 594 => b"00000_0000_00_001010010111", -- load, gr0, YPOS2
 595 => b"00011_0000_01_000000000000", -- sub, gr0
 596 => b"00000_0000_00_000000000001", -- 1
 597 => b"01000_0000_01_000000000000", -- mul, gr0
 598 => b"00000_0000_00_000000001111", -- 15
 599 => b"00010_0000_00_001010010110", -- add, gr0, XPOS2
 600 => b"10000_0000_00_000000000000", -- tpoint, gr0
 601 => b"01111_0001_00_000000000000", -- tread, gr1
 602 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 603 => b"00111_0000_01_000000000000", -- bne
 604 => b"00000_0000_00_000000000100", -- CONTROL_R
 605 => b"00011_1111_01_000000000000", -- sub, gr15
 606 => b"00000_0000_00_000000000001", -- 1
 607 => b"00100_0000_01_000000000000", -- jump
 608 => b"00000_0000_00_000000000100", -- CONTROL_R
 609 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 610 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 611 => b"00000_0000_00_001010010111", -- load, gr0, YPOS2
 612 => b"01000_0000_01_000000000000", -- mul, gr0
 613 => b"00000_0000_00_000000001111", -- 15
 614 => b"00010_0000_00_001010010110", -- add, gr0, XPOS2
 615 => b"00011_0000_01_000000000000", -- sub, gr0
 616 => b"00000_0000_00_000000000001", -- 1
 617 => b"10000_0000_00_000000000000", -- tpoint, gr0
 618 => b"01111_0001_00_000000000000", -- tread, gr1
 619 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 620 => b"00111_0000_01_000000000000", -- bne
 621 => b"00000_0000_00_000111110101", -- J3
 622 => b"00011_1110_01_000000000000", -- sub, gr14
 623 => b"00000_0000_00_000000000001", -- 1
 624 => b"00100_0000_01_000000000000", -- jump
 625 => b"00000_0000_00_000111110101", -- J3
 626 => b"00001_1110_10_001010010110", -- store, gr14, XPOS2
 627 => b"00001_1111_10_001010010111", -- store, gr15, YPOS2
 628 => b"00000_0000_00_001010010111", -- load, gr0, YPOS2
 629 => b"00010_0000_01_000000000000", -- add, gr0
 630 => b"00000_0000_00_000000000001", -- 1
 631 => b"01000_0000_01_000000000000", -- mul, gr0
 632 => b"00000_0000_00_000000001111", -- 15
 633 => b"00010_0000_00_001010010110", -- add, gr0, XPOS2
 634 => b"10000_0000_00_000000000000", -- tpoint, gr0
 635 => b"01111_0001_00_000000000000", -- tread, gr1
 636 => b"00011_0001_00_001010011011", -- sub, gr1, GRASS
 637 => b"00111_0000_01_000000000000", -- bne
 638 => b"00000_0000_00_000000000100", -- CONTROL_R
 639 => b"00010_1111_01_000000000000", -- add, gr15
 640 => b"00000_0000_00_000000000001", -- 1
 641 => b"00100_0000_01_000000000000", -- jump
 642 => b"00000_0000_00_000000000100", -- CONTROL_R
 643 => b"00100_0000_01_000000000000", -- jump
 644 => b"00000_0000_00_000111101001", -- COUNT_R
 645 => b"00000_0000_00_000000000000", -- 0
 646 => b"00000_0000_00_000000000000", -- 0
 647 => b"00000_0000_00_000000000000", -- 0
 648 => b"00000_0000_00_000000000000", -- 0
 649 => b"00000_0000_00_000000000000", -- 0
 650 => b"00000_0000_00_000000000000", -- 0
 651 => b"00000_0000_00_000000000000", -- 0
 652 => b"00000_0000_00_000000000000", -- 0
 653 => b"00000_0000_00_000000000000", -- 0
 654 => b"00000_0000_00_000000000000", -- 0
 655 => b"00000_0000_00_000000000000", -- 0
 656 => b"00000_0000_00_000000000000", -- 0
 657 => b"00000_0000_00_000000000000", -- 0
 658 => b"00000_0000_00_000000000000", -- 0
 659 => b"00000_0000_00_000000000001", -- 1
 660 => b"00000_0000_00_000000000000", -- 0
 661 => b"00000_0000_00_000000000000", -- 0
 662 => b"00000_0000_00_000000000000", -- 0
 663 => b"00000_0000_00_000000000000", -- 0
 664 => b"00000_0000_00_000000000000", -- 0
 665 => b"00000_0000_00_000000000000", -- 0
 666 => b"00000_0000_00_000000000000", -- 0
 667 => b"00000_0000_00_000000000000", -- 0
 668 => b"00000_0000_00_000000000001", -- 1
 669 => b"00000_0000_00_000000000010", -- 2
 670 => b"00000_0000_00_000000000011", -- 3
 671 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
