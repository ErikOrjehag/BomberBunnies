library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_001010010001", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000111010101", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011000100", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000010000", -- BOOM1
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000001101010", -- BOOM2
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  16 => b"00000_0000_00_001100110011", -- load, gr0, P1EXPLOSION1ACTIVE
  17 => b"00011_0000_01_000000000000", -- sub, gr0
  18 => b"00000_0000_00_000000000001", -- 1
  19 => b"00111_0000_01_000000000000", -- bne
  20 => b"00000_0000_00_000000001100", -- BOOM1_R
  21 => b"00000_0000_00_001100110010", -- load, gr0, P1EXPLOSION1TIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000001", -- 1
  24 => b"00001_0000_10_001100110010", -- store, gr0, P1EXPLOSION1TIME
  25 => b"00000_0000_00_001100110010", -- load, gr0, P1EXPLOSION1TIME
  26 => b"00011_0000_01_000000000000", -- sub, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00111_0000_01_000000000000", -- bne
  29 => b"00000_0000_00_000000001100", -- BOOM1_R
  30 => b"00000_0000_01_000000000000", -- load, gr0
  31 => b"00000_0000_00_000000000000", -- 0
  32 => b"00001_0000_10_001100110011", -- store, gr0, P1EXPLOSION1ACTIVE
  33 => b"00000_0010_00_001100110100", -- load, gr2, P1EXPLOSION1POS
  34 => b"00000_0011_00_001101011101", -- load, gr3, GRASS
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01110_0011_00_000000000000", -- twrite, gr3
  37 => b"00010_0010_01_000000000000", -- add, gr2
  38 => b"00000_0000_00_000000000001", -- 1
  39 => b"10000_0010_00_000000000000", -- tpoint, gr2
  40 => b"01111_0000_00_000000000000", -- tread, gr0
  41 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  42 => b"00111_0000_01_000000000000", -- bne
  43 => b"00000_0000_00_000000110101", -- E1LEFT
  44 => b"01110_0011_00_000000000000", -- twrite, gr3
  45 => b"00010_0010_01_000000000000", -- add, gr2
  46 => b"00000_0000_00_000000000001", -- 1
  47 => b"10000_0010_00_000000000000", -- tpoint, gr2
  48 => b"01111_0000_00_000000000000", -- tread, gr0
  49 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  50 => b"00111_0000_01_000000000000", -- bne
  51 => b"00000_0000_00_000000110101", -- E1LEFT
  52 => b"01110_0011_00_000000000000", -- twrite, gr3
  53 => b"00000_0010_00_001100110100", -- load, gr2, P1EXPLOSION1POS
  54 => b"00011_0010_01_000000000000", -- sub, gr2
  55 => b"00000_0000_00_000000000001", -- 1
  56 => b"10000_0010_00_000000000000", -- tpoint, gr2
  57 => b"01111_0000_00_000000000000", -- tread, gr0
  58 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  59 => b"00111_0000_01_000000000000", -- bne
  60 => b"00000_0000_00_000001000110", -- E1DOWN
  61 => b"01110_0011_00_000000000000", -- twrite, gr3
  62 => b"00011_0010_01_000000000000", -- sub, gr2
  63 => b"00000_0000_00_000000000001", -- 1
  64 => b"10000_0010_00_000000000000", -- tpoint, gr2
  65 => b"01111_0000_00_000000000000", -- tread, gr0
  66 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  67 => b"00111_0000_01_000000000000", -- bne
  68 => b"00000_0000_00_000001000110", -- E1DOWN
  69 => b"01110_0011_00_000000000000", -- twrite, gr3
  70 => b"00000_0010_00_001100110100", -- load, gr2, P1EXPLOSION1POS
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000001111", -- 15
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0000_00_000000000000", -- tread, gr0
  75 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  76 => b"00111_0000_01_000000000000", -- bne
  77 => b"00000_0000_00_000001010111", -- E1UP
  78 => b"01110_0011_00_000000000000", -- twrite, gr3
  79 => b"00010_0010_01_000000000000", -- add, gr2
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"10000_0010_00_000000000000", -- tpoint, gr2
  82 => b"01111_0000_00_000000000000", -- tread, gr0
  83 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  84 => b"00111_0000_01_000000000000", -- bne
  85 => b"00000_0000_00_000001010111", -- E1UP
  86 => b"01110_0011_00_000000000000", -- twrite, gr3
  87 => b"00000_0010_00_001100110100", -- load, gr2, P1EXPLOSION1POS
  88 => b"00011_0010_01_000000000000", -- sub, gr2
  89 => b"00000_0000_00_000000001111", -- 15
  90 => b"10000_0010_00_000000000000", -- tpoint, gr2
  91 => b"01111_0000_00_000000000000", -- tread, gr0
  92 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
  93 => b"00111_0000_01_000000000000", -- bne
  94 => b"00000_0000_00_000000001100", -- BOOM1_R
  95 => b"01110_0011_00_000000000000", -- twrite, gr3
  96 => b"00011_0010_01_000000000000", -- sub, gr2
  97 => b"00000_0000_00_000000001111", -- 15
  98 => b"10000_0010_00_000000000000", -- tpoint, gr2
  99 => b"01111_0000_00_000000000000", -- tread, gr0
 100 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 101 => b"00111_0000_01_000000000000", -- bne
 102 => b"00000_0000_00_000000001100", -- BOOM1_R
 103 => b"01110_0011_00_000000000000", -- twrite, gr3
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000000001100", -- BOOM1_R
 106 => b"00000_0000_00_001101000101", -- load, gr0, P2EXPLOSION1ACTIVE
 107 => b"00011_0000_01_000000000000", -- sub, gr0
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00111_0000_01_000000000000", -- bne
 110 => b"00000_0000_00_000000001110", -- BOOM2_R
 111 => b"00000_0000_00_001101000100", -- load, gr0, P2EXPLOSION1TIME
 112 => b"00011_0000_01_000000000000", -- sub, gr0
 113 => b"00000_0000_00_000000000001", -- 1
 114 => b"00001_0000_10_001101000100", -- store, gr0, P2EXPLOSION1TIME
 115 => b"00000_0000_00_001101000100", -- load, gr0, P2EXPLOSION1TIME
 116 => b"00011_0000_01_000000000000", -- sub, gr0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00111_0000_01_000000000000", -- bne
 119 => b"00000_0000_00_000000001110", -- BOOM2_R
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001101000101", -- store, gr0, P2EXPLOSION1ACTIVE
 123 => b"00000_0010_00_001101000110", -- load, gr2, P2EXPLOSION1POS
 124 => b"00000_0011_00_001101011101", -- load, gr3, GRASS
 125 => b"10000_0010_00_000000000000", -- tpoint, gr2
 126 => b"01110_0011_00_000000000000", -- twrite, gr3
 127 => b"00010_0010_01_000000000000", -- add, gr2
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"10000_0010_00_000000000000", -- tpoint, gr2
 130 => b"01111_0000_00_000000000000", -- tread, gr0
 131 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 132 => b"00111_0000_01_000000000000", -- bne
 133 => b"00000_0000_00_000010001111", -- E2LEFT
 134 => b"01110_0011_00_000000000000", -- twrite, gr3
 135 => b"00010_0010_01_000000000000", -- add, gr2
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0010_00_000000000000", -- tpoint, gr2
 138 => b"01111_0000_00_000000000000", -- tread, gr0
 139 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000010001111", -- E2LEFT
 142 => b"01110_0011_00_000000000000", -- twrite, gr3
 143 => b"00000_0010_00_001101000110", -- load, gr2, P2EXPLOSION1POS
 144 => b"00011_0010_01_000000000000", -- sub, gr2
 145 => b"00000_0000_00_000000000001", -- 1
 146 => b"10000_0010_00_000000000000", -- tpoint, gr2
 147 => b"01111_0000_00_000000000000", -- tread, gr0
 148 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 149 => b"00111_0000_01_000000000000", -- bne
 150 => b"00000_0000_00_000010100000", -- E2DOWN
 151 => b"01110_0011_00_000000000000", -- twrite, gr3
 152 => b"00011_0010_01_000000000000", -- sub, gr2
 153 => b"00000_0000_00_000000000001", -- 1
 154 => b"10000_0010_00_000000000000", -- tpoint, gr2
 155 => b"01111_0000_00_000000000000", -- tread, gr0
 156 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000010100000", -- E2DOWN
 159 => b"01110_0011_00_000000000000", -- twrite, gr3
 160 => b"00000_0010_00_001101000110", -- load, gr2, P2EXPLOSION1POS
 161 => b"00010_0010_01_000000000000", -- add, gr2
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"10000_0010_00_000000000000", -- tpoint, gr2
 164 => b"01111_0000_00_000000000000", -- tread, gr0
 165 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 166 => b"00111_0000_01_000000000000", -- bne
 167 => b"00000_0000_00_000010110001", -- E2UP
 168 => b"01110_0011_00_000000000000", -- twrite, gr3
 169 => b"00010_0010_01_000000000000", -- add, gr2
 170 => b"00000_0000_00_000000001111", -- 15
 171 => b"10000_0010_00_000000000000", -- tpoint, gr2
 172 => b"01111_0000_00_000000000000", -- tread, gr0
 173 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000010110001", -- E2UP
 176 => b"01110_0011_00_000000000000", -- twrite, gr3
 177 => b"00000_0010_00_001101000110", -- load, gr2, P2EXPLOSION1POS
 178 => b"00011_0010_01_000000000000", -- sub, gr2
 179 => b"00000_0000_00_000000001111", -- 15
 180 => b"10000_0010_00_000000000000", -- tpoint, gr2
 181 => b"01111_0000_00_000000000000", -- tread, gr0
 182 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 183 => b"00111_0000_01_000000000000", -- bne
 184 => b"00000_0000_00_000000001110", -- BOOM2_R
 185 => b"01110_0011_00_000000000000", -- twrite, gr3
 186 => b"00011_0010_01_000000000000", -- sub, gr2
 187 => b"00000_0000_00_000000001111", -- 15
 188 => b"10000_0010_00_000000000000", -- tpoint, gr2
 189 => b"01111_0000_00_000000000000", -- tread, gr0
 190 => b"00011_0000_00_001101100000", -- sub, gr0, EXPLOSION
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000001110", -- BOOM2_R
 193 => b"01110_0011_00_000000000000", -- twrite, gr3
 194 => b"00100_0000_01_000000000000", -- jump
 195 => b"00000_0000_00_000000001110", -- BOOM2_R
 196 => b"00000_0000_00_001100110001", -- load, gr0, P1BOMB1ACTIVE
 197 => b"00011_0000_01_000000000000", -- sub, gr0
 198 => b"00000_0000_00_000000000001", -- 1
 199 => b"00111_0000_01_000000000000", -- bne
 200 => b"00000_0000_00_000011010010", -- P1BOMB2
 201 => b"00000_0000_00_001100110000", -- load, gr0, P1BOMB1TIME
 202 => b"00011_0000_01_000000000000", -- sub, gr0
 203 => b"00000_0000_00_000000000001", -- 1
 204 => b"00001_0000_10_001100110000", -- store, gr0, P1BOMB1TIME
 205 => b"00000_0000_01_000000000000", -- load, gr0
 206 => b"00000_0000_00_000000000000", -- 0
 207 => b"00011_0000_00_001100110000", -- sub, gr0, P1BOMB1TIME
 208 => b"00110_0000_01_000000000000", -- beq
 209 => b"00000_0000_00_000100011100", -- P1EXPLOSION1INIT
 210 => b"00000_0000_00_001100110111", -- load, gr0, P1BOMB2ACTIVE
 211 => b"00011_0000_01_000000000000", -- sub, gr0
 212 => b"00000_0000_00_000000000001", -- 1
 213 => b"00111_0000_01_000000000000", -- bne
 214 => b"00000_0000_00_000011100000", -- P1BOMB3
 215 => b"00000_0000_00_001100110110", -- load, gr0, P1BOMB2TIME
 216 => b"00011_0000_01_000000000000", -- sub, gr0
 217 => b"00000_0000_00_000000000001", -- 1
 218 => b"00001_0000_10_001100110110", -- store, gr0, P1BOMB2TIME
 219 => b"00000_0000_01_000000000000", -- load, gr0
 220 => b"00000_0000_00_000000000000", -- 0
 221 => b"00011_0000_00_001100110110", -- sub, gr0, P1BOMB2TIME
 222 => b"00110_0000_01_000000000000", -- beq
 223 => b"00000_0000_00_000100101110", -- P1EXPLOSION2INIT
 224 => b"00000_0000_00_001100111101", -- load, gr0, P1BOMB3ACTIVE
 225 => b"00011_0000_01_000000000000", -- sub, gr0
 226 => b"00000_0000_00_000000000001", -- 1
 227 => b"00111_0000_01_000000000000", -- bne
 228 => b"00000_0000_00_000011110000", -- P2BOMB1
 229 => b"00000_0000_00_001100111100", -- load, gr0, P1BOMB3TIME
 230 => b"00011_0000_01_000000000000", -- sub, gr0
 231 => b"00000_0000_00_000000000001", -- 1
 232 => b"00001_0000_10_001100111100", -- store, gr0, P1BOMB3TIME
 233 => b"00000_0000_01_000000000000", -- load, gr0
 234 => b"00000_0000_00_000000000000", -- 0
 235 => b"00011_0000_00_001100111100", -- sub, gr0, P1BOMB3TIME
 236 => b"00110_0000_01_000000000000", -- beq
 237 => b"00000_0000_00_000101000000", -- P1EXPLOSION3INIT
 238 => b"00100_0000_01_000000000000", -- jump
 239 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 240 => b"00000_0000_00_001101000011", -- load, gr0, P2BOMB1ACTIVE
 241 => b"00011_0000_01_000000000000", -- sub, gr0
 242 => b"00000_0000_00_000000000001", -- 1
 243 => b"00111_0000_01_000000000000", -- bne
 244 => b"00000_0000_00_000011111110", -- P2BOMB2
 245 => b"00000_0000_00_001101000010", -- load, gr0, P2BOMB1TIME
 246 => b"00011_0000_01_000000000000", -- sub, gr0
 247 => b"00000_0000_00_000000000001", -- 1
 248 => b"00001_0000_10_001101000010", -- store, gr0, P2BOMB1TIME
 249 => b"00000_0000_01_000000000000", -- load, gr0
 250 => b"00000_0000_00_000000000000", -- 0
 251 => b"00011_0000_00_001101000010", -- sub, gr0, P2BOMB1TIME
 252 => b"00110_0000_01_000000000000", -- beq
 253 => b"00000_0000_00_000101010010", -- P2EXPLOSION1INIT
 254 => b"00000_0000_00_001101001001", -- load, gr0, P2BOMB2ACTIVE
 255 => b"00011_0000_01_000000000000", -- sub, gr0
 256 => b"00000_0000_00_000000000001", -- 1
 257 => b"00111_0000_01_000000000000", -- bne
 258 => b"00000_0000_00_000100001100", -- P2BOMB3
 259 => b"00000_0000_00_001101001000", -- load, gr0, P2BOMB2TIME
 260 => b"00011_0000_01_000000000000", -- sub, gr0
 261 => b"00000_0000_00_000000000001", -- 1
 262 => b"00001_0000_10_001101001000", -- store, gr0, P2BOMB2TIME
 263 => b"00000_0000_01_000000000000", -- load, gr0
 264 => b"00000_0000_00_000000000000", -- 0
 265 => b"00011_0000_00_001101001000", -- sub, gr0, P2BOMB2TIME
 266 => b"00110_0000_01_000000000000", -- beq
 267 => b"00000_0000_00_000101100100", -- P2EXPLOSION2INIT
 268 => b"00000_0000_00_001101001111", -- load, gr0, P2BOMB3ACTIVE
 269 => b"00011_0000_01_000000000000", -- sub, gr0
 270 => b"00000_0000_00_000000000001", -- 1
 271 => b"00111_0000_01_000000000000", -- bne
 272 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 273 => b"00000_0000_00_001101001110", -- load, gr0, P2BOMB3TIME
 274 => b"00011_0000_01_000000000000", -- sub, gr0
 275 => b"00000_0000_00_000000000001", -- 1
 276 => b"00001_0000_10_001101001110", -- store, gr0, P2BOMB3TIME
 277 => b"00000_0000_01_000000000000", -- load, gr0
 278 => b"00000_0000_00_000000000000", -- 0
 279 => b"00011_0000_00_001101001110", -- sub, gr0, P2BOMB3TIME
 280 => b"00110_0000_01_000000000000", -- beq
 281 => b"00000_0000_00_000101110110", -- P2EXPLOSION3INIT
 282 => b"00100_0000_01_000000000000", -- jump
 283 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 284 => b"00000_0000_01_000000000000", -- load, gr0
 285 => b"00000_0000_00_000000000000", -- 0
 286 => b"00001_0000_10_001100110001", -- store, gr0, P1BOMB1ACTIVE
 287 => b"00000_0000_00_001100101111", -- load, gr0, P1BOMB1POS
 288 => b"00001_0000_10_001100110100", -- store, gr0, P1EXPLOSION1POS
 289 => b"00000_0000_01_000000000000", -- load, gr0
 290 => b"00000_0000_00_000000000001", -- 1
 291 => b"00001_0000_10_001100110011", -- store, gr0, P1EXPLOSION1ACTIVE
 292 => b"00000_0000_01_000000000000", -- load, gr0
 293 => b"00000_0000_00_000000000010", -- 2
 294 => b"00001_0000_10_001100110010", -- store, gr0, P1EXPLOSION1TIME
 295 => b"00000_0000_00_001101010011", -- load, gr0, P1BOMBCOUNT
 296 => b"00011_0000_01_000000000000", -- sub, gr0
 297 => b"00000_0000_00_000000000001", -- 1
 298 => b"00001_0000_10_001101010011", -- store, gr0, P1BOMBCOUNT
 299 => b"00000_0100_00_001100101111", -- load, gr4, P1BOMB1POS
 300 => b"00100_0000_01_000000000000", -- jump
 301 => b"00000_0000_00_000110001000", -- EXPLODE
 302 => b"00000_0000_01_000000000000", -- load, gr0
 303 => b"00000_0000_00_000000000000", -- 0
 304 => b"00001_0000_10_001100110111", -- store, gr0, P1BOMB2ACTIVE
 305 => b"00000_0000_00_001100110101", -- load, gr0, P1BOMB2POS
 306 => b"00001_0000_10_001100111010", -- store, gr0, P1EXPLOSION2POS
 307 => b"00000_0000_01_000000000000", -- load, gr0
 308 => b"00000_0000_00_000000000001", -- 1
 309 => b"00001_0000_10_001100111001", -- store, gr0, P1EXPLOSION2ACTIVE
 310 => b"00000_0000_01_000000000000", -- load, gr0
 311 => b"00000_0000_00_000000000010", -- 2
 312 => b"00001_0000_10_001100111000", -- store, gr0, P1EXPLOSION2TIME
 313 => b"00000_0000_00_001101010011", -- load, gr0, P1BOMBCOUNT
 314 => b"00011_0000_01_000000000000", -- sub, gr0
 315 => b"00000_0000_00_000000000001", -- 1
 316 => b"00001_0000_10_001101010011", -- store, gr0, P1BOMBCOUNT
 317 => b"00000_0100_00_001100110101", -- load, gr4, P1BOMB2POS
 318 => b"00100_0000_01_000000000000", -- jump
 319 => b"00000_0000_00_000110001000", -- EXPLODE
 320 => b"00000_0000_01_000000000000", -- load, gr0
 321 => b"00000_0000_00_000000000000", -- 0
 322 => b"00001_0000_10_001100111101", -- store, gr0, P1BOMB3ACTIVE
 323 => b"00000_0000_00_001100111011", -- load, gr0, P1BOMB3POS
 324 => b"00001_0000_10_001101000000", -- store, gr0, P1EXPLOSION3POS
 325 => b"00000_0000_01_000000000000", -- load, gr0
 326 => b"00000_0000_00_000000000001", -- 1
 327 => b"00001_0000_10_001100111111", -- store, gr0, P1EXPLOSION3ACTIVE
 328 => b"00000_0000_01_000000000000", -- load, gr0
 329 => b"00000_0000_00_000000000010", -- 2
 330 => b"00001_0000_10_001100111110", -- store, gr0, P1EXPLOSION3TIME
 331 => b"00000_0000_00_001101010011", -- load, gr0, P1BOMBCOUNT
 332 => b"00011_0000_01_000000000000", -- sub, gr0
 333 => b"00000_0000_00_000000000001", -- 1
 334 => b"00001_0000_10_001101010011", -- store, gr0, P1BOMBCOUNT
 335 => b"00000_0100_00_001100111011", -- load, gr4, P1BOMB3POS
 336 => b"00100_0000_01_000000000000", -- jump
 337 => b"00000_0000_00_000110001000", -- EXPLODE
 338 => b"00000_0000_01_000000000000", -- load, gr0
 339 => b"00000_0000_00_000000000000", -- 0
 340 => b"00001_0000_10_001101000011", -- store, gr0, P2BOMB1ACTIVE
 341 => b"00000_0000_00_001101000001", -- load, gr0, P2BOMB1POS
 342 => b"00001_0000_10_001101000110", -- store, gr0, P2EXPLOSION1POS
 343 => b"00000_0000_01_000000000000", -- load, gr0
 344 => b"00000_0000_00_000000000001", -- 1
 345 => b"00001_0000_10_001101000101", -- store, gr0, P2EXPLOSION1ACTIVE
 346 => b"00000_0000_01_000000000000", -- load, gr0
 347 => b"00000_0000_00_000000000010", -- 2
 348 => b"00001_0000_10_001101000100", -- store, gr0, P2EXPLOSION1TIME
 349 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMBCOUNT
 350 => b"00011_0000_01_000000000000", -- sub, gr0
 351 => b"00000_0000_00_000000000001", -- 1
 352 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMBCOUNT
 353 => b"00000_0100_00_001101000001", -- load, gr4, P2BOMB1POS
 354 => b"00100_0000_01_000000000000", -- jump
 355 => b"00000_0000_00_000110001000", -- EXPLODE
 356 => b"00000_0000_01_000000000000", -- load, gr0
 357 => b"00000_0000_00_000000000000", -- 0
 358 => b"00001_0000_10_001101001001", -- store, gr0, P2BOMB2ACTIVE
 359 => b"00000_0000_00_001101000111", -- load, gr0, P2BOMB2POS
 360 => b"00001_0000_10_001101001100", -- store, gr0, P2EXPLOSION2POS
 361 => b"00000_0000_01_000000000000", -- load, gr0
 362 => b"00000_0000_00_000000000001", -- 1
 363 => b"00001_0000_10_001101001011", -- store, gr0, P2EXPLOSION2ACTIVE
 364 => b"00000_0000_01_000000000000", -- load, gr0
 365 => b"00000_0000_00_000000000010", -- 2
 366 => b"00001_0000_10_001101001010", -- store, gr0, P2EXPLOSION2TIME
 367 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMBCOUNT
 368 => b"00011_0000_01_000000000000", -- sub, gr0
 369 => b"00000_0000_00_000000000001", -- 1
 370 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMBCOUNT
 371 => b"00000_0100_00_001101000111", -- load, gr4, P2BOMB2POS
 372 => b"00100_0000_01_000000000000", -- jump
 373 => b"00000_0000_00_000110001000", -- EXPLODE
 374 => b"00000_0000_01_000000000000", -- load, gr0
 375 => b"00000_0000_00_000000000000", -- 0
 376 => b"00001_0000_10_001101001111", -- store, gr0, P2BOMB3ACTIVE
 377 => b"00000_0000_00_001101001101", -- load, gr0, P2BOMB3POS
 378 => b"00001_0000_10_001101010010", -- store, gr0, P2EXPLOSION3POS
 379 => b"00000_0000_01_000000000000", -- load, gr0
 380 => b"00000_0000_00_000000000001", -- 1
 381 => b"00001_0000_10_001101010001", -- store, gr0, P2EXPLOSION3ACTIVE
 382 => b"00000_0000_01_000000000000", -- load, gr0
 383 => b"00000_0000_00_000000000010", -- 2
 384 => b"00001_0000_10_001101010000", -- store, gr0, P2EXPLOSION3TIME
 385 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMBCOUNT
 386 => b"00011_0000_01_000000000000", -- sub, gr0
 387 => b"00000_0000_00_000000000001", -- 1
 388 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMBCOUNT
 389 => b"00000_0100_00_001101001101", -- load, gr4, P2BOMB3POS
 390 => b"00100_0000_01_000000000000", -- jump
 391 => b"00000_0000_00_000110001000", -- EXPLODE
 392 => b"00001_0100_10_001101011010", -- store, gr4, MOVE
 393 => b"00000_0010_00_001101011010", -- load, gr2, MOVE
 394 => b"00000_0011_00_001101100000", -- load, gr3, EXPLOSION
 395 => b"10000_0010_00_000000000000", -- tpoint, gr2
 396 => b"01110_0011_00_000000000000", -- twrite, gr3
 397 => b"00010_0010_01_000000000000", -- add, gr2
 398 => b"00000_0000_00_000000000001", -- 1
 399 => b"10000_0010_00_000000000000", -- tpoint, gr2
 400 => b"01111_0000_00_000000000000", -- tread, gr0
 401 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 402 => b"00110_0000_01_000000000000", -- beq
 403 => b"00000_0000_00_000110011101", -- EXPLODELEFT
 404 => b"01110_0011_00_000000000000", -- twrite, gr3
 405 => b"00010_0010_01_000000000000", -- add, gr2
 406 => b"00000_0000_00_000000000001", -- 1
 407 => b"10000_0010_00_000000000000", -- tpoint, gr2
 408 => b"01111_0000_00_000000000000", -- tread, gr0
 409 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 410 => b"00110_0000_01_000000000000", -- beq
 411 => b"00000_0000_00_000110011101", -- EXPLODELEFT
 412 => b"01110_0011_00_000000000000", -- twrite, gr3
 413 => b"00001_0100_10_001101011010", -- store, gr4, MOVE
 414 => b"00000_0010_00_001101011010", -- load, gr2, MOVE
 415 => b"00011_0010_01_000000000000", -- sub, gr2
 416 => b"00000_0000_00_000000000001", -- 1
 417 => b"10000_0010_00_000000000000", -- tpoint, gr2
 418 => b"01111_0000_00_000000000000", -- tread, gr0
 419 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 420 => b"00110_0000_01_000000000000", -- beq
 421 => b"00000_0000_00_000110101111", -- EXPLODEDOWN
 422 => b"01110_0011_00_000000000000", -- twrite, gr3
 423 => b"00011_0010_01_000000000000", -- sub, gr2
 424 => b"00000_0000_00_000000000001", -- 1
 425 => b"10000_0010_00_000000000000", -- tpoint, gr2
 426 => b"01111_0000_00_000000000000", -- tread, gr0
 427 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 428 => b"00110_0000_01_000000000000", -- beq
 429 => b"00000_0000_00_000110101111", -- EXPLODEDOWN
 430 => b"01110_0011_00_000000000000", -- twrite, gr3
 431 => b"00001_0100_10_001101011010", -- store, gr4, MOVE
 432 => b"00000_0010_00_001101011010", -- load, gr2, MOVE
 433 => b"00010_0010_01_000000000000", -- add, gr2
 434 => b"00000_0000_00_000000001111", -- 15
 435 => b"10000_0010_00_000000000000", -- tpoint, gr2
 436 => b"01111_0000_00_000000000000", -- tread, gr0
 437 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 438 => b"00110_0000_01_000000000000", -- beq
 439 => b"00000_0000_00_000111000001", -- EXPLODEUP
 440 => b"01110_0011_00_000000000000", -- twrite, gr3
 441 => b"00010_0010_01_000000000000", -- add, gr2
 442 => b"00000_0000_00_000000001111", -- 15
 443 => b"10000_0010_00_000000000000", -- tpoint, gr2
 444 => b"01111_0000_00_000000000000", -- tread, gr0
 445 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 446 => b"00110_0000_01_000000000000", -- beq
 447 => b"00000_0000_00_000111000001", -- EXPLODEUP
 448 => b"01110_0011_00_000000000000", -- twrite, gr3
 449 => b"00001_0100_10_001101011010", -- store, gr4, MOVE
 450 => b"00000_0010_00_001101011010", -- load, gr2, MOVE
 451 => b"00011_0010_01_000000000000", -- sub, gr2
 452 => b"00000_0000_00_000000001111", -- 15
 453 => b"10000_0010_00_000000000000", -- tpoint, gr2
 454 => b"01111_0000_00_000000000000", -- tread, gr0
 455 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 456 => b"00110_0000_01_000000000000", -- beq
 457 => b"00000_0000_00_000011000100", -- TICKBOMBS
 458 => b"01110_0011_00_000000000000", -- twrite, gr3
 459 => b"00011_0010_01_000000000000", -- sub, gr2
 460 => b"00000_0000_00_000000001111", -- 15
 461 => b"10000_0010_00_000000000000", -- tpoint, gr2
 462 => b"01111_0000_00_000000000000", -- tread, gr0
 463 => b"00011_0000_00_001101011110", -- sub, gr0, WALL
 464 => b"00110_0000_01_000000000000", -- beq
 465 => b"00000_0000_00_000011000100", -- TICKBOMBS
 466 => b"01110_0011_00_000000000000", -- twrite, gr3
 467 => b"00100_0000_01_000000000000", -- jump
 468 => b"00000_0000_00_000011000100", -- TICKBOMBS
 469 => b"10101_0000_01_000000000000", -- btn1
 470 => b"00000_0000_00_000111011011", -- BTN1
 471 => b"11010_0000_01_000000000000", -- btn2
 472 => b"00000_0000_00_001000110111", -- BTN2
 473 => b"00100_0000_01_000000000000", -- jump
 474 => b"00000_0000_00_000000000100", -- BUTTON_R
 475 => b"00000_0000_00_001101010011", -- load, gr0, P1BOMBCOUNT
 476 => b"00011_0000_00_001101010101", -- sub, gr0, MAXBOMBS
 477 => b"00110_0000_01_000000000000", -- beq
 478 => b"00000_0000_00_000111010111", -- BTN1_R
 479 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 480 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 481 => b"00000_0000_00_001101010111", -- load, gr0, YPOS1
 482 => b"01000_0000_01_000000000000", -- mul, gr0
 483 => b"00000_0000_00_000000001111", -- 15
 484 => b"00010_0000_00_001101010110", -- add, gr0, XPOS1
 485 => b"10000_0000_00_000000000000", -- tpoint, gr0
 486 => b"01111_0001_00_000000000000", -- tread, gr1
 487 => b"00011_0001_00_001101100001", -- sub, gr1, EGG
 488 => b"00110_0000_01_000000000000", -- beq
 489 => b"00000_0000_00_000111010111", -- BTN1_R
 490 => b"00000_0000_00_001100110001", -- load, gr0, P1BOMB1ACTIVE
 491 => b"00011_0000_01_000000000000", -- sub, gr0
 492 => b"00000_0000_00_000000000000", -- 0
 493 => b"00110_0000_01_000000000000", -- beq
 494 => b"00000_0000_00_001000000001", -- P1PLACEBOMB1
 495 => b"00000_0000_00_001100110111", -- load, gr0, P1BOMB2ACTIVE
 496 => b"00011_0000_01_000000000000", -- sub, gr0
 497 => b"00000_0000_00_000000000000", -- 0
 498 => b"00110_0000_01_000000000000", -- beq
 499 => b"00000_0000_00_001000010011", -- P1PLACEBOMB2
 500 => b"00000_0000_00_001100111101", -- load, gr0, P1BOMB3ACTIVE
 501 => b"00011_0000_01_000000000000", -- sub, gr0
 502 => b"00000_0000_00_000000000000", -- 0
 503 => b"00110_0000_01_000000000000", -- beq
 504 => b"00000_0000_00_001000100101", -- P1PLACEBOMB3
 505 => b"00100_0000_01_000000000000", -- jump
 506 => b"00000_0000_00_000111010111", -- BTN1_R
 507 => b"00000_0000_00_001101010011", -- load, gr0, P1BOMBCOUNT
 508 => b"00010_0000_01_000000000000", -- add, gr0
 509 => b"00000_0000_00_000000000001", -- 1
 510 => b"00001_0000_10_001101010011", -- store, gr0, P1BOMBCOUNT
 511 => b"00100_0000_01_000000000000", -- jump
 512 => b"00000_0000_00_000111010111", -- BTN1_R
 513 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 514 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 515 => b"00000_0011_00_001101010111", -- load, gr3, YPOS1
 516 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 517 => b"01000_0011_01_000000000000", -- mul, gr3
 518 => b"00000_0000_00_000000001111", -- 15
 519 => b"00010_0011_00_001101010110", -- add, gr3, XPOS1
 520 => b"10000_0011_00_000000000000", -- tpoint, gr3
 521 => b"01110_0010_00_000000000000", -- twrite, gr2
 522 => b"00000_0000_01_000000000000", -- load, gr0
 523 => b"00000_0000_00_000000000001", -- 1
 524 => b"00001_0000_10_001100110001", -- store, gr0, P1BOMB1ACTIVE
 525 => b"00001_0011_10_001100101111", -- store, gr3, P1BOMB1POS
 526 => b"00000_0000_01_000000000000", -- load, gr0
 527 => b"00000_0000_00_000000010000", -- 16
 528 => b"00001_0000_10_001100110000", -- store, gr0, P1BOMB1TIME
 529 => b"00100_0000_01_000000000000", -- jump
 530 => b"00000_0000_00_000111111011", -- P1INCREASEBOMBCOUNTER
 531 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 532 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 533 => b"00000_0011_00_001101010111", -- load, gr3, YPOS1
 534 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 535 => b"01000_0011_01_000000000000", -- mul, gr3
 536 => b"00000_0000_00_000000001111", -- 15
 537 => b"00010_0011_00_001101010110", -- add, gr3, XPOS1
 538 => b"10000_0011_00_000000000000", -- tpoint, gr3
 539 => b"01110_0010_00_000000000000", -- twrite, gr2
 540 => b"00000_0000_01_000000000000", -- load, gr0
 541 => b"00000_0000_00_000000000001", -- 1
 542 => b"00001_0000_10_001100110111", -- store, gr0, P1BOMB2ACTIVE
 543 => b"00001_0011_10_001100110101", -- store, gr3, P1BOMB2POS
 544 => b"00000_0000_01_000000000000", -- load, gr0
 545 => b"00000_0000_00_000000010000", -- 16
 546 => b"00001_0000_10_001100110110", -- store, gr0, P1BOMB2TIME
 547 => b"00100_0000_01_000000000000", -- jump
 548 => b"00000_0000_00_000111111011", -- P1INCREASEBOMBCOUNTER
 549 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 550 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 551 => b"00000_0011_00_001101010111", -- load, gr3, YPOS1
 552 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 553 => b"01000_0011_01_000000000000", -- mul, gr3
 554 => b"00000_0000_00_000000001111", -- 15
 555 => b"00010_0011_00_001101010110", -- add, gr3, XPOS1
 556 => b"10000_0011_00_000000000000", -- tpoint, gr3
 557 => b"01110_0010_00_000000000000", -- twrite, gr2
 558 => b"00000_0000_01_000000000000", -- load, gr0
 559 => b"00000_0000_00_000000000001", -- 1
 560 => b"00001_0000_10_001100111101", -- store, gr0, P1BOMB3ACTIVE
 561 => b"00001_0011_10_001100111011", -- store, gr3, P1BOMB3POS
 562 => b"00000_0000_01_000000000000", -- load, gr0
 563 => b"00000_0000_00_000000010000", -- 16
 564 => b"00001_0000_10_001100111100", -- store, gr0, P1BOMB3TIME
 565 => b"00100_0000_01_000000000000", -- jump
 566 => b"00000_0000_00_000111111011", -- P1INCREASEBOMBCOUNTER
 567 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMBCOUNT
 568 => b"00011_0000_00_001101010101", -- sub, gr0, MAXBOMBS
 569 => b"00110_0000_01_000000000000", -- beq
 570 => b"00000_0000_00_000111011001", -- BTN2_R
 571 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 572 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 573 => b"00000_0000_00_001101011001", -- load, gr0, YPOS2
 574 => b"01000_0000_01_000000000000", -- mul, gr0
 575 => b"00000_0000_00_000000001111", -- 15
 576 => b"00010_0000_00_001101011000", -- add, gr0, XPOS2
 577 => b"10000_0000_00_000000000000", -- tpoint, gr0
 578 => b"01111_0001_00_000000000000", -- tread, gr1
 579 => b"00011_0001_00_001101100001", -- sub, gr1, EGG
 580 => b"00110_0000_01_000000000000", -- beq
 581 => b"00000_0000_00_000111011001", -- BTN2_R
 582 => b"00000_0000_00_001101000011", -- load, gr0, P2BOMB1ACTIVE
 583 => b"00011_0000_01_000000000000", -- sub, gr0
 584 => b"00000_0000_00_000000000000", -- 0
 585 => b"00110_0000_01_000000000000", -- beq
 586 => b"00000_0000_00_001001011011", -- P2PLACEBOMB1
 587 => b"00000_0000_00_001101001001", -- load, gr0, P2BOMB2ACTIVE
 588 => b"00011_0000_01_000000000000", -- sub, gr0
 589 => b"00000_0000_00_000000000000", -- 0
 590 => b"00110_0000_01_000000000000", -- beq
 591 => b"00000_0000_00_001001101101", -- P2PLACEBOMB2
 592 => b"00000_0000_00_001101001111", -- load, gr0, P2BOMB3ACTIVE
 593 => b"00011_0000_01_000000000000", -- sub, gr0
 594 => b"00000_0000_00_000000000000", -- 0
 595 => b"00110_0000_01_000000000000", -- beq
 596 => b"00000_0000_00_001001111111", -- P2PLACEBOMB3
 597 => b"00000_0000_00_001101010100", -- load, gr0, P2BOMBCOUNT
 598 => b"00010_0000_01_000000000000", -- add, gr0
 599 => b"00000_0000_00_000000000001", -- 1
 600 => b"00001_0000_10_001101010100", -- store, gr0, P2BOMBCOUNT
 601 => b"00100_0000_01_000000000000", -- jump
 602 => b"00000_0000_00_000111011001", -- BTN2_R
 603 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 604 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 605 => b"00000_0011_00_001101011001", -- load, gr3, YPOS2
 606 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 607 => b"01000_0011_01_000000000000", -- mul, gr3
 608 => b"00000_0000_00_000000001111", -- 15
 609 => b"00010_0011_00_001101011000", -- add, gr3, XPOS2
 610 => b"10000_0011_00_000000000000", -- tpoint, gr3
 611 => b"01110_0010_00_000000000000", -- twrite, gr2
 612 => b"00000_0000_01_000000000000", -- load, gr0
 613 => b"00000_0000_00_000000000001", -- 1
 614 => b"00001_0000_10_001101000011", -- store, gr0, P2BOMB1ACTIVE
 615 => b"00001_0011_10_001101000001", -- store, gr3, P2BOMB1POS
 616 => b"00000_0000_01_000000000000", -- load, gr0
 617 => b"00000_0000_00_000000010000", -- 16
 618 => b"00001_0000_10_001101000010", -- store, gr0, P2BOMB1TIME
 619 => b"00100_0000_01_000000000000", -- jump
 620 => b"00000_0000_00_001001010101", -- P2INCREASEBOMBCOUNTER
 621 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 622 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 623 => b"00000_0011_00_001101011001", -- load, gr3, YPOS2
 624 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 625 => b"01000_0011_01_000000000000", -- mul, gr3
 626 => b"00000_0000_00_000000001111", -- 15
 627 => b"00010_0011_00_001101011000", -- add, gr3, XPOS2
 628 => b"10000_0011_00_000000000000", -- tpoint, gr3
 629 => b"01110_0010_00_000000000000", -- twrite, gr2
 630 => b"00000_0000_01_000000000000", -- load, gr0
 631 => b"00000_0000_00_000000000001", -- 1
 632 => b"00001_0000_10_001101001001", -- store, gr0, P2BOMB2ACTIVE
 633 => b"00001_0011_10_001101000111", -- store, gr3, P2BOMB2POS
 634 => b"00000_0000_01_000000000000", -- load, gr0
 635 => b"00000_0000_00_000000010000", -- 16
 636 => b"00001_0000_10_001101001000", -- store, gr0, P2BOMB2TIME
 637 => b"00100_0000_01_000000000000", -- jump
 638 => b"00000_0000_00_001001010101", -- P2INCREASEBOMBCOUNTER
 639 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 640 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 641 => b"00000_0011_00_001101011001", -- load, gr3, YPOS2
 642 => b"00000_0010_00_001101100001", -- load, gr2, EGG
 643 => b"01000_0011_01_000000000000", -- mul, gr3
 644 => b"00000_0000_00_000000001111", -- 15
 645 => b"00010_0011_00_001101011000", -- add, gr3, XPOS2
 646 => b"10000_0011_00_000000000000", -- tpoint, gr3
 647 => b"01110_0010_00_000000000000", -- twrite, gr2
 648 => b"00000_0000_01_000000000000", -- load, gr0
 649 => b"00000_0000_00_000000000001", -- 1
 650 => b"00001_0000_10_001101001111", -- store, gr0, P2BOMB3ACTIVE
 651 => b"00001_0011_10_001101001101", -- store, gr3, P2BOMB3POS
 652 => b"00000_0000_01_000000000000", -- load, gr0
 653 => b"00000_0000_00_000000010000", -- 16
 654 => b"00001_0000_10_001101001110", -- store, gr0, P2BOMB3TIME
 655 => b"00100_0000_01_000000000000", -- jump
 656 => b"00000_0000_00_001001010101", -- P2INCREASEBOMBCOUNTER
 657 => b"00100_0000_01_000000000000", -- jump
 658 => b"00000_0000_00_001100101101", -- COUNT1
 659 => b"10001_0000_01_000000000000", -- joy1r
 660 => b"00000_0000_00_001010100101", -- P1R
 661 => b"10011_0000_01_000000000000", -- joy1l
 662 => b"00000_0000_00_001011000111", -- P1L
 663 => b"10010_0000_01_000000000000", -- joy1u
 664 => b"00000_0000_00_001010110110", -- P1U
 665 => b"10100_0000_01_000000000000", -- joy1d
 666 => b"00000_0000_00_001011011000", -- P1D
 667 => b"10110_0000_01_000000000000", -- joy2r
 668 => b"00000_0000_00_001011101001", -- P2R
 669 => b"11000_0000_01_000000000000", -- joy2l
 670 => b"00000_0000_00_001100001011", -- P2L
 671 => b"10111_0000_01_000000000000", -- joy2u
 672 => b"00000_0000_00_001011111010", -- P2U
 673 => b"11001_0000_01_000000000000", -- joy2d
 674 => b"00000_0000_00_001100011100", -- P2D
 675 => b"00100_0000_01_000000000000", -- jump
 676 => b"00000_0000_00_000000000010", -- CONTROL_R
 677 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 678 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 679 => b"00000_0000_00_001101010111", -- load, gr0, YPOS1
 680 => b"01000_0000_01_000000000000", -- mul, gr0
 681 => b"00000_0000_00_000000001111", -- 15
 682 => b"00010_0000_00_001101010110", -- add, gr0, XPOS1
 683 => b"00010_0000_01_000000000000", -- add, gr0
 684 => b"00000_0000_00_000000000001", -- 1
 685 => b"10000_0000_00_000000000000", -- tpoint, gr0
 686 => b"01111_0001_00_000000000000", -- tread, gr1
 687 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 688 => b"00111_0000_01_000000000000", -- bne
 689 => b"00000_0000_00_001010010111", -- J1
 690 => b"00010_1100_01_000000000000", -- add, gr12
 691 => b"00000_0000_00_000000000001", -- 1
 692 => b"00100_0000_01_000000000000", -- jump
 693 => b"00000_0000_00_001010010111", -- J1
 694 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 695 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 696 => b"00000_0000_00_001101010111", -- load, gr0, YPOS1
 697 => b"00011_0000_01_000000000000", -- sub, gr0
 698 => b"00000_0000_00_000000000001", -- 1
 699 => b"01000_0000_01_000000000000", -- mul, gr0
 700 => b"00000_0000_00_000000001111", -- 15
 701 => b"00010_0000_00_001101010110", -- add, gr0, XPOS1
 702 => b"10000_0000_00_000000000000", -- tpoint, gr0
 703 => b"01111_0001_00_000000000000", -- tread, gr1
 704 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 705 => b"00111_0000_01_000000000000", -- bne
 706 => b"00000_0000_00_001010011011", -- J2
 707 => b"00011_1101_01_000000000000", -- sub, gr13
 708 => b"00000_0000_00_000000000001", -- 1
 709 => b"00100_0000_01_000000000000", -- jump
 710 => b"00000_0000_00_001010011011", -- J2
 711 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 712 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 713 => b"00000_0000_00_001101010111", -- load, gr0, YPOS1
 714 => b"01000_0000_01_000000000000", -- mul, gr0
 715 => b"00000_0000_00_000000001111", -- 15
 716 => b"00010_0000_00_001101010110", -- add, gr0, XPOS1
 717 => b"00011_0000_01_000000000000", -- sub, gr0
 718 => b"00000_0000_00_000000000001", -- 1
 719 => b"10000_0000_00_000000000000", -- tpoint, gr0
 720 => b"01111_0001_00_000000000000", -- tread, gr1
 721 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 722 => b"00111_0000_01_000000000000", -- bne
 723 => b"00000_0000_00_001010010111", -- J1
 724 => b"00011_1100_01_000000000000", -- sub, gr12
 725 => b"00000_0000_00_000000000001", -- 1
 726 => b"00100_0000_01_000000000000", -- jump
 727 => b"00000_0000_00_001010010111", -- J1
 728 => b"00001_1100_10_001101010110", -- store, gr12, XPOS1
 729 => b"00001_1101_10_001101010111", -- store, gr13, YPOS1
 730 => b"00000_0000_00_001101010111", -- load, gr0, YPOS1
 731 => b"00010_0000_01_000000000000", -- add, gr0
 732 => b"00000_0000_00_000000000001", -- 1
 733 => b"01000_0000_01_000000000000", -- mul, gr0
 734 => b"00000_0000_00_000000001111", -- 15
 735 => b"00010_0000_00_001101010110", -- add, gr0, XPOS1
 736 => b"10000_0000_00_000000000000", -- tpoint, gr0
 737 => b"01111_0001_00_000000000000", -- tread, gr1
 738 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 739 => b"00111_0000_01_000000000000", -- bne
 740 => b"00000_0000_00_001010011011", -- J2
 741 => b"00010_1101_01_000000000000", -- add, gr13
 742 => b"00000_0000_00_000000000001", -- 1
 743 => b"00100_0000_01_000000000000", -- jump
 744 => b"00000_0000_00_001010011011", -- J2
 745 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 746 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 747 => b"00000_0000_00_001101011001", -- load, gr0, YPOS2
 748 => b"01000_0000_01_000000000000", -- mul, gr0
 749 => b"00000_0000_00_000000001111", -- 15
 750 => b"00010_0000_00_001101011000", -- add, gr0, XPOS2
 751 => b"00010_0000_01_000000000000", -- add, gr0
 752 => b"00000_0000_00_000000000001", -- 1
 753 => b"10000_0000_00_000000000000", -- tpoint, gr0
 754 => b"01111_0001_00_000000000000", -- tread, gr1
 755 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 756 => b"00111_0000_01_000000000000", -- bne
 757 => b"00000_0000_00_001010011111", -- J3
 758 => b"00010_1110_01_000000000000", -- add, gr14
 759 => b"00000_0000_00_000000000001", -- 1
 760 => b"00100_0000_01_000000000000", -- jump
 761 => b"00000_0000_00_001010011111", -- J3
 762 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 763 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 764 => b"00000_0000_00_001101011001", -- load, gr0, YPOS2
 765 => b"00011_0000_01_000000000000", -- sub, gr0
 766 => b"00000_0000_00_000000000001", -- 1
 767 => b"01000_0000_01_000000000000", -- mul, gr0
 768 => b"00000_0000_00_000000001111", -- 15
 769 => b"00010_0000_00_001101011000", -- add, gr0, XPOS2
 770 => b"10000_0000_00_000000000000", -- tpoint, gr0
 771 => b"01111_0001_00_000000000000", -- tread, gr1
 772 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 773 => b"00111_0000_01_000000000000", -- bne
 774 => b"00000_0000_00_000000000010", -- CONTROL_R
 775 => b"00011_1111_01_000000000000", -- sub, gr15
 776 => b"00000_0000_00_000000000001", -- 1
 777 => b"00100_0000_01_000000000000", -- jump
 778 => b"00000_0000_00_000000000010", -- CONTROL_R
 779 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 780 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 781 => b"00000_0000_00_001101011001", -- load, gr0, YPOS2
 782 => b"01000_0000_01_000000000000", -- mul, gr0
 783 => b"00000_0000_00_000000001111", -- 15
 784 => b"00010_0000_00_001101011000", -- add, gr0, XPOS2
 785 => b"00011_0000_01_000000000000", -- sub, gr0
 786 => b"00000_0000_00_000000000001", -- 1
 787 => b"10000_0000_00_000000000000", -- tpoint, gr0
 788 => b"01111_0001_00_000000000000", -- tread, gr1
 789 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 790 => b"00111_0000_01_000000000000", -- bne
 791 => b"00000_0000_00_001010011111", -- J3
 792 => b"00011_1110_01_000000000000", -- sub, gr14
 793 => b"00000_0000_00_000000000001", -- 1
 794 => b"00100_0000_01_000000000000", -- jump
 795 => b"00000_0000_00_001010011111", -- J3
 796 => b"00001_1110_10_001101011000", -- store, gr14, XPOS2
 797 => b"00001_1111_10_001101011001", -- store, gr15, YPOS2
 798 => b"00000_0000_00_001101011001", -- load, gr0, YPOS2
 799 => b"00010_0000_01_000000000000", -- add, gr0
 800 => b"00000_0000_00_000000000001", -- 1
 801 => b"01000_0000_01_000000000000", -- mul, gr0
 802 => b"00000_0000_00_000000001111", -- 15
 803 => b"00010_0000_00_001101011000", -- add, gr0, XPOS2
 804 => b"10000_0000_00_000000000000", -- tpoint, gr0
 805 => b"01111_0001_00_000000000000", -- tread, gr1
 806 => b"00011_0001_00_001101011101", -- sub, gr1, GRASS
 807 => b"00111_0000_01_000000000000", -- bne
 808 => b"00000_0000_00_000000000010", -- CONTROL_R
 809 => b"00010_1111_01_000000000000", -- add, gr15
 810 => b"00000_0000_00_000000000001", -- 1
 811 => b"00100_0000_01_000000000000", -- jump
 812 => b"00000_0000_00_000000000010", -- CONTROL_R
 813 => b"00100_0000_01_000000000000", -- jump
 814 => b"00000_0000_00_001010010011", -- COUNT_R
 815 => b"00000_0000_00_000000000000", -- 0
 816 => b"00000_0000_00_000000000000", -- 0
 817 => b"00000_0000_00_000000000000", -- 0
 818 => b"00000_0000_00_000000000000", -- 0
 819 => b"00000_0000_00_000000000000", -- 0
 820 => b"00000_0000_00_000000000000", -- 0
 821 => b"00000_0000_00_000000000000", -- 0
 822 => b"00000_0000_00_000000000000", -- 0
 823 => b"00000_0000_00_000000000000", -- 0
 824 => b"00000_0000_00_000000000000", -- 0
 825 => b"00000_0000_00_000000000000", -- 0
 826 => b"00000_0000_00_000000000000", -- 0
 827 => b"00000_0000_00_000000000000", -- 0
 828 => b"00000_0000_00_000000000000", -- 0
 829 => b"00000_0000_00_000000000000", -- 0
 830 => b"00000_0000_00_000000000000", -- 0
 831 => b"00000_0000_00_000000000000", -- 0
 832 => b"00000_0000_00_000000000000", -- 0
 833 => b"00000_0000_00_000000000000", -- 0
 834 => b"00000_0000_00_000000000000", -- 0
 835 => b"00000_0000_00_000000000000", -- 0
 836 => b"00000_0000_00_000000000000", -- 0
 837 => b"00000_0000_00_000000000000", -- 0
 838 => b"00000_0000_00_000000000000", -- 0
 839 => b"00000_0000_00_000000000000", -- 0
 840 => b"00000_0000_00_000000000000", -- 0
 841 => b"00000_0000_00_000000000000", -- 0
 842 => b"00000_0000_00_000000000000", -- 0
 843 => b"00000_0000_00_000000000000", -- 0
 844 => b"00000_0000_00_000000000000", -- 0
 845 => b"00000_0000_00_000000000000", -- 0
 846 => b"00000_0000_00_000000000000", -- 0
 847 => b"00000_0000_00_000000000000", -- 0
 848 => b"00000_0000_00_000000000000", -- 0
 849 => b"00000_0000_00_000000000000", -- 0
 850 => b"00000_0000_00_000000000000", -- 0
 851 => b"00000_0000_00_000000000000", -- 0
 852 => b"00000_0000_00_000000000000", -- 0
 853 => b"00000_0000_00_000000000011", -- 3
 854 => b"00000_0000_00_000000000000", -- 0
 855 => b"00000_0000_00_000000000000", -- 0
 856 => b"00000_0000_00_000000000000", -- 0
 857 => b"00000_0000_00_000000000000", -- 0
 858 => b"00000_0000_00_000000000000", -- 0
 859 => b"00000_0000_00_000000000000", -- 0
 860 => b"00000_0000_00_000000000000", -- 0
 861 => b"00000_0000_00_000000000000", -- 0
 862 => b"00000_0000_00_000000000001", -- 1
 863 => b"00000_0000_00_000000000010", -- 2
 864 => b"00000_0000_00_000000000011", -- 3
 865 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
