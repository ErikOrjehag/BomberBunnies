library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000100", -- 4
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000110000111", -- CONTROL
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000100110110", -- BUTTON
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000001100110", -- TICKBOMBS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000001100", -- TICKEXPLOSIONS
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000000010", -- MAIN
  12 => b"00000_0000_00_001000101001", -- load, gr0, P1EXPLOSIONACTIVE
  13 => b"00011_0000_01_000000000000", -- sub, gr0
  14 => b"00000_0000_00_000000000001", -- 1
  15 => b"00111_0000_01_000000000000", -- bne
  16 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  17 => b"00000_0000_00_001000101000", -- load, gr0, P1EXPLOSIONTIME
  18 => b"00011_0000_01_000000000000", -- sub, gr0
  19 => b"00000_0000_00_000000000001", -- 1
  20 => b"00001_0000_10_001000101000", -- store, gr0, P1EXPLOSIONTIME
  21 => b"00000_0000_00_001000101000", -- load, gr0, P1EXPLOSIONTIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000000", -- 0
  24 => b"00111_0000_01_000000000000", -- bne
  25 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  26 => b"00000_0000_01_000000000000", -- load, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00001_0000_10_001000101001", -- store, gr0, P1EXPLOSIONACTIVE
  29 => b"00000_0010_00_001000101010", -- load, gr2, P1EXPLOSIONPOS
  30 => b"00000_0011_00_001000111011", -- load, gr3, GRASS
  31 => b"10000_0010_00_000000000000", -- tpoint, gr2
  32 => b"01110_0011_00_000000000000", -- twrite, gr3
  33 => b"00010_0010_01_000000000000", -- add, gr2
  34 => b"00000_0000_00_000000000001", -- 1
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01111_0000_00_000000000000", -- tread, gr0
  37 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  38 => b"00111_0000_01_000000000000", -- bne
  39 => b"00000_0000_00_000000110001", -- E1LEFT
  40 => b"01110_0011_00_000000000000", -- twrite, gr3
  41 => b"00010_0010_01_000000000000", -- add, gr2
  42 => b"00000_0000_00_000000000001", -- 1
  43 => b"10000_0010_00_000000000000", -- tpoint, gr2
  44 => b"01111_0000_00_000000000000", -- tread, gr0
  45 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  46 => b"00111_0000_01_000000000000", -- bne
  47 => b"00000_0000_00_000000110001", -- E1LEFT
  48 => b"01110_0011_00_000000000000", -- twrite, gr3
  49 => b"00000_0010_00_001000101010", -- load, gr2, P1EXPLOSIONPOS
  50 => b"00011_0010_01_000000000000", -- sub, gr2
  51 => b"00000_0000_00_000000000001", -- 1
  52 => b"10000_0010_00_000000000000", -- tpoint, gr2
  53 => b"01111_0000_00_000000000000", -- tread, gr0
  54 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  55 => b"00111_0000_01_000000000000", -- bne
  56 => b"00000_0000_00_000001000010", -- E1DOWN
  57 => b"01110_0011_00_000000000000", -- twrite, gr3
  58 => b"00011_0010_01_000000000000", -- sub, gr2
  59 => b"00000_0000_00_000000000001", -- 1
  60 => b"10000_0010_00_000000000000", -- tpoint, gr2
  61 => b"01111_0000_00_000000000000", -- tread, gr0
  62 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  63 => b"00111_0000_01_000000000000", -- bne
  64 => b"00000_0000_00_000001000010", -- E1DOWN
  65 => b"01110_0011_00_000000000000", -- twrite, gr3
  66 => b"00000_0010_00_001000101010", -- load, gr2, P1EXPLOSIONPOS
  67 => b"00010_0010_01_000000000000", -- add, gr2
  68 => b"00000_0000_00_000000001111", -- 15
  69 => b"10000_0010_00_000000000000", -- tpoint, gr2
  70 => b"01111_0000_00_000000000000", -- tread, gr0
  71 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  72 => b"00111_0000_01_000000000000", -- bne
  73 => b"00000_0000_00_000001010011", -- E1UP
  74 => b"01110_0011_00_000000000000", -- twrite, gr3
  75 => b"00010_0010_01_000000000000", -- add, gr2
  76 => b"00000_0000_00_000000001111", -- 15
  77 => b"10000_0010_00_000000000000", -- tpoint, gr2
  78 => b"01111_0000_00_000000000000", -- tread, gr0
  79 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  80 => b"00111_0000_01_000000000000", -- bne
  81 => b"00000_0000_00_000001010011", -- E1UP
  82 => b"01110_0011_00_000000000000", -- twrite, gr3
  83 => b"00000_0010_00_001000101010", -- load, gr2, P1EXPLOSIONPOS
  84 => b"00011_0010_01_000000000000", -- sub, gr2
  85 => b"00000_0000_00_000000001111", -- 15
  86 => b"10000_0010_00_000000000000", -- tpoint, gr2
  87 => b"01111_0000_00_000000000000", -- tread, gr0
  88 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  89 => b"00111_0000_01_000000000000", -- bne
  90 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  91 => b"01110_0011_00_000000000000", -- twrite, gr3
  92 => b"00011_0010_01_000000000000", -- sub, gr2
  93 => b"00000_0000_00_000000001111", -- 15
  94 => b"10000_0010_00_000000000000", -- tpoint, gr2
  95 => b"01111_0000_00_000000000000", -- tread, gr0
  96 => b"00011_0000_00_001000111110", -- sub, gr0, EXPLOSION
  97 => b"00111_0000_01_000000000000", -- bne
  98 => b"00000_0000_00_000001100100", -- TICKEXPLOSION2
  99 => b"01110_0011_00_000000000000", -- twrite, gr3
 100 => b"00100_0000_01_000000000000", -- jump
 101 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS_R
 102 => b"00100_0000_01_000000000000", -- jump
 103 => b"00000_0000_00_000001101100", -- TICKBOMB1
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000011010001", -- TICKBOMB2
 106 => b"00100_0000_01_000000000000", -- jump
 107 => b"00000_0000_00_000000001000", -- TICKBOMBS_R
 108 => b"00000_0000_00_001000100111", -- load, gr0, P1BOMBACTIVE
 109 => b"00011_0000_01_000000000000", -- sub, gr0
 110 => b"00000_0000_00_000000000001", -- 1
 111 => b"00111_0000_01_000000000000", -- bne
 112 => b"00000_0000_00_000001101000", -- TICKBOMB1_R
 113 => b"00000_0000_00_001000100110", -- load, gr0, P1BOMBTIME
 114 => b"00011_0000_01_000000000000", -- sub, gr0
 115 => b"00000_0000_00_000000000001", -- 1
 116 => b"00001_0000_10_001000100110", -- store, gr0, P1BOMBTIME
 117 => b"00000_0000_01_000000000000", -- load, gr0
 118 => b"00000_0000_00_000000000000", -- 0
 119 => b"00011_0000_00_001000100110", -- sub, gr0, P1BOMBTIME
 120 => b"00110_0000_01_000000000000", -- beq
 121 => b"00000_0000_00_000001111100", -- EXPLODE1
 122 => b"00100_0000_01_000000000000", -- jump
 123 => b"00000_0000_00_000001101000", -- TICKBOMB1_R
 124 => b"00000_0000_00_001000100101", -- load, gr0, P1BOMBPOS
 125 => b"00001_0000_10_001000101010", -- store, gr0, P1EXPLOSIONPOS
 126 => b"00000_0000_01_000000000000", -- load, gr0
 127 => b"00000_0000_00_000000000001", -- 1
 128 => b"00001_0000_10_001000101001", -- store, gr0, P1EXPLOSIONACTIVE
 129 => b"00000_0000_01_000000000000", -- load, gr0
 130 => b"00000_0000_00_000000000010", -- 2
 131 => b"00001_0000_10_001000101000", -- store, gr0, P1EXPLOSIONTIME
 132 => b"00000_0000_00_001000110001", -- load, gr0, BOMBS1
 133 => b"00011_0000_01_000000000000", -- sub, gr0
 134 => b"00000_0000_00_000000000001", -- 1
 135 => b"00001_0000_10_001000110001", -- store, gr0, BOMBS1
 136 => b"00000_0010_00_001000100101", -- load, gr2, P1BOMBPOS
 137 => b"00000_0011_00_001000111110", -- load, gr3, EXPLOSION
 138 => b"10000_0010_00_000000000000", -- tpoint, gr2
 139 => b"01110_0011_00_000000000000", -- twrite, gr3
 140 => b"00010_0010_01_000000000000", -- add, gr2
 141 => b"00000_0000_00_000000000001", -- 1
 142 => b"10000_0010_00_000000000000", -- tpoint, gr2
 143 => b"01111_0000_00_000000000000", -- tread, gr0
 144 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 145 => b"00110_0000_01_000000000000", -- beq
 146 => b"00000_0000_00_000010011100", -- P1LEFT
 147 => b"01110_0011_00_000000000000", -- twrite, gr3
 148 => b"00010_0010_01_000000000000", -- add, gr2
 149 => b"00000_0000_00_000000000001", -- 1
 150 => b"10000_0010_00_000000000000", -- tpoint, gr2
 151 => b"01111_0000_00_000000000000", -- tread, gr0
 152 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 153 => b"00110_0000_01_000000000000", -- beq
 154 => b"00000_0000_00_000010011100", -- P1LEFT
 155 => b"01110_0011_00_000000000000", -- twrite, gr3
 156 => b"00000_0010_00_001000100101", -- load, gr2, P1BOMBPOS
 157 => b"00011_0010_01_000000000000", -- sub, gr2
 158 => b"00000_0000_00_000000000001", -- 1
 159 => b"10000_0010_00_000000000000", -- tpoint, gr2
 160 => b"01111_0000_00_000000000000", -- tread, gr0
 161 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 162 => b"00110_0000_01_000000000000", -- beq
 163 => b"00000_0000_00_000010101101", -- P1DOWN
 164 => b"01110_0011_00_000000000000", -- twrite, gr3
 165 => b"00011_0010_01_000000000000", -- sub, gr2
 166 => b"00000_0000_00_000000000001", -- 1
 167 => b"10000_0010_00_000000000000", -- tpoint, gr2
 168 => b"01111_0000_00_000000000000", -- tread, gr0
 169 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 170 => b"00110_0000_01_000000000000", -- beq
 171 => b"00000_0000_00_000010101101", -- P1DOWN
 172 => b"01110_0011_00_000000000000", -- twrite, gr3
 173 => b"00000_0010_00_001000100101", -- load, gr2, P1BOMBPOS
 174 => b"00010_0010_01_000000000000", -- add, gr2
 175 => b"00000_0000_00_000000001111", -- 15
 176 => b"10000_0010_00_000000000000", -- tpoint, gr2
 177 => b"01111_0000_00_000000000000", -- tread, gr0
 178 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 179 => b"00110_0000_01_000000000000", -- beq
 180 => b"00000_0000_00_000010111110", -- P1UP
 181 => b"01110_0011_00_000000000000", -- twrite, gr3
 182 => b"00010_0010_01_000000000000", -- add, gr2
 183 => b"00000_0000_00_000000001111", -- 15
 184 => b"10000_0010_00_000000000000", -- tpoint, gr2
 185 => b"01111_0000_00_000000000000", -- tread, gr0
 186 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 187 => b"00110_0000_01_000000000000", -- beq
 188 => b"00000_0000_00_000010111110", -- P1UP
 189 => b"01110_0011_00_000000000000", -- twrite, gr3
 190 => b"00000_0010_00_001000100101", -- load, gr2, P1BOMBPOS
 191 => b"00011_0010_01_000000000000", -- sub, gr2
 192 => b"00000_0000_00_000000001111", -- 15
 193 => b"10000_0010_00_000000000000", -- tpoint, gr2
 194 => b"01111_0000_00_000000000000", -- tread, gr0
 195 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 196 => b"00110_0000_01_000000000000", -- beq
 197 => b"00000_0000_00_000001101000", -- TICKBOMB1_R
 198 => b"01110_0011_00_000000000000", -- twrite, gr3
 199 => b"00011_0010_01_000000000000", -- sub, gr2
 200 => b"00000_0000_00_000000001111", -- 15
 201 => b"10000_0010_00_000000000000", -- tpoint, gr2
 202 => b"01111_0000_00_000000000000", -- tread, gr0
 203 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 204 => b"00110_0000_01_000000000000", -- beq
 205 => b"00000_0000_00_000001101000", -- TICKBOMB1_R
 206 => b"01110_0011_00_000000000000", -- twrite, gr3
 207 => b"00100_0000_01_000000000000", -- jump
 208 => b"00000_0000_00_000001101000", -- TICKBOMB1_R
 209 => b"00000_0000_00_001000101101", -- load, gr0, P2BOMBACTIVE
 210 => b"00011_0000_01_000000000000", -- sub, gr0
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00111_0000_01_000000000000", -- bne
 213 => b"00000_0000_00_000001101010", -- TICKBOMB2_R
 214 => b"00000_0000_00_001000101100", -- load, gr0, P2BOMBTIME
 215 => b"00011_0000_01_000000000000", -- sub, gr0
 216 => b"00000_0000_00_000000000001", -- 1
 217 => b"00001_0000_10_001000101100", -- store, gr0, P2BOMBTIME
 218 => b"00000_0000_01_000000000000", -- load, gr0
 219 => b"00000_0000_00_000000000000", -- 0
 220 => b"00011_0000_00_001000101100", -- sub, gr0, P2BOMBTIME
 221 => b"00110_0000_01_000000000000", -- beq
 222 => b"00000_0000_00_000011100001", -- EXPLODE2
 223 => b"00100_0000_01_000000000000", -- jump
 224 => b"00000_0000_00_000001101010", -- TICKBOMB2_R
 225 => b"00000_0000_00_001000101011", -- load, gr0, P2BOMBPOS
 226 => b"00001_0000_10_001000110000", -- store, gr0, P2EXPLOSIONPOS
 227 => b"00000_0000_01_000000000000", -- load, gr0
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00001_0000_10_001000101111", -- store, gr0, P2EXPLOSIONACTIVE
 230 => b"00000_0000_01_000000000000", -- load, gr0
 231 => b"00000_0000_00_000000000010", -- 2
 232 => b"00001_0000_10_001000101110", -- store, gr0, P2EXPLOSIONTIME
 233 => b"00000_0000_00_001000110010", -- load, gr0, BOMBS2
 234 => b"00011_0000_01_000000000000", -- sub, gr0
 235 => b"00000_0000_00_000000000001", -- 1
 236 => b"00001_0000_10_001000110010", -- store, gr0, BOMBS2
 237 => b"00000_0010_00_001000101011", -- load, gr2, P2BOMBPOS
 238 => b"00000_0011_00_001000111110", -- load, gr3, EXPLOSION
 239 => b"10000_0010_00_000000000000", -- tpoint, gr2
 240 => b"01110_0011_00_000000000000", -- twrite, gr3
 241 => b"00010_0010_01_000000000000", -- add, gr2
 242 => b"00000_0000_00_000000000001", -- 1
 243 => b"10000_0010_00_000000000000", -- tpoint, gr2
 244 => b"01111_0000_00_000000000000", -- tread, gr0
 245 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 246 => b"00110_0000_01_000000000000", -- beq
 247 => b"00000_0000_00_000100000001", -- P2LEFT
 248 => b"01110_0011_00_000000000000", -- twrite, gr3
 249 => b"00010_0010_01_000000000000", -- add, gr2
 250 => b"00000_0000_00_000000000001", -- 1
 251 => b"10000_0010_00_000000000000", -- tpoint, gr2
 252 => b"01111_0000_00_000000000000", -- tread, gr0
 253 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 254 => b"00110_0000_01_000000000000", -- beq
 255 => b"00000_0000_00_000100000001", -- P2LEFT
 256 => b"01110_0011_00_000000000000", -- twrite, gr3
 257 => b"00000_0010_00_001000101011", -- load, gr2, P2BOMBPOS
 258 => b"00011_0010_01_000000000000", -- sub, gr2
 259 => b"00000_0000_00_000000000001", -- 1
 260 => b"10000_0010_00_000000000000", -- tpoint, gr2
 261 => b"01111_0000_00_000000000000", -- tread, gr0
 262 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 263 => b"00110_0000_01_000000000000", -- beq
 264 => b"00000_0000_00_000100010010", -- P2DOWN
 265 => b"01110_0011_00_000000000000", -- twrite, gr3
 266 => b"00011_0010_01_000000000000", -- sub, gr2
 267 => b"00000_0000_00_000000000001", -- 1
 268 => b"10000_0010_00_000000000000", -- tpoint, gr2
 269 => b"01111_0000_00_000000000000", -- tread, gr0
 270 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 271 => b"00110_0000_01_000000000000", -- beq
 272 => b"00000_0000_00_000100010010", -- P2DOWN
 273 => b"01110_0011_00_000000000000", -- twrite, gr3
 274 => b"00000_0010_00_001000101011", -- load, gr2, P2BOMBPOS
 275 => b"00010_0010_01_000000000000", -- add, gr2
 276 => b"00000_0000_00_000000001111", -- 15
 277 => b"10000_0010_00_000000000000", -- tpoint, gr2
 278 => b"01111_0000_00_000000000000", -- tread, gr0
 279 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 280 => b"00110_0000_01_000000000000", -- beq
 281 => b"00000_0000_00_000100100011", -- P2UP
 282 => b"01110_0011_00_000000000000", -- twrite, gr3
 283 => b"00010_0010_01_000000000000", -- add, gr2
 284 => b"00000_0000_00_000000001111", -- 15
 285 => b"10000_0010_00_000000000000", -- tpoint, gr2
 286 => b"01111_0000_00_000000000000", -- tread, gr0
 287 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 288 => b"00110_0000_01_000000000000", -- beq
 289 => b"00000_0000_00_000100100011", -- P2UP
 290 => b"01110_0011_00_000000000000", -- twrite, gr3
 291 => b"00000_0010_00_001000101011", -- load, gr2, P2BOMBPOS
 292 => b"00011_0010_01_000000000000", -- sub, gr2
 293 => b"00000_0000_00_000000001111", -- 15
 294 => b"10000_0010_00_000000000000", -- tpoint, gr2
 295 => b"01111_0000_00_000000000000", -- tread, gr0
 296 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 297 => b"00110_0000_01_000000000000", -- beq
 298 => b"00000_0000_00_000001101010", -- TICKBOMB2_R
 299 => b"01110_0011_00_000000000000", -- twrite, gr3
 300 => b"00011_0010_01_000000000000", -- sub, gr2
 301 => b"00000_0000_00_000000001111", -- 15
 302 => b"10000_0010_00_000000000000", -- tpoint, gr2
 303 => b"01111_0000_00_000000000000", -- tread, gr0
 304 => b"00011_0000_00_001000111100", -- sub, gr0, WALL
 305 => b"00110_0000_01_000000000000", -- beq
 306 => b"00000_0000_00_000001101010", -- TICKBOMB2_R
 307 => b"01110_0011_00_000000000000", -- twrite, gr3
 308 => b"00100_0000_01_000000000000", -- jump
 309 => b"00000_0000_00_000001101010", -- TICKBOMB2_R
 310 => b"10101_0000_01_000000000000", -- btn1
 311 => b"00000_0000_00_000100111100", -- BTN1
 312 => b"11010_0000_01_000000000000", -- btn2
 313 => b"00000_0000_00_000101100001", -- BTN2
 314 => b"00100_0000_01_000000000000", -- jump
 315 => b"00000_0000_00_000000000110", -- BUTTON_R
 316 => b"00000_0000_00_001000110001", -- load, gr0, BOMBS1
 317 => b"00011_0000_00_001000110011", -- sub, gr0, MAXBOMBS
 318 => b"00110_0000_01_000000000000", -- beq
 319 => b"00000_0000_00_000100111000", -- BTN1_R
 320 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 321 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 322 => b"00000_0000_00_001000110101", -- load, gr0, YPOS1
 323 => b"01000_0000_01_000000000000", -- mul, gr0
 324 => b"00000_0000_00_000000001111", -- 15
 325 => b"00010_0000_00_001000110100", -- add, gr0, XPOS1
 326 => b"10000_0000_00_000000000000", -- tpoint, gr0
 327 => b"01111_0001_00_000000000000", -- tread, gr1
 328 => b"00011_0001_00_001000111111", -- sub, gr1, EGG
 329 => b"00110_0000_01_000000000000", -- beq
 330 => b"00000_0000_00_000100111000", -- BTN1_R
 331 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 332 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 333 => b"00000_0011_00_001000110101", -- load, gr3, YPOS1
 334 => b"00000_0010_00_001000111111", -- load, gr2, EGG
 335 => b"01000_0011_01_000000000000", -- mul, gr3
 336 => b"00000_0000_00_000000001111", -- 15
 337 => b"00010_0011_00_001000110100", -- add, gr3, XPOS1
 338 => b"10000_0011_00_000000000000", -- tpoint, gr3
 339 => b"01110_0010_00_000000000000", -- twrite, gr2
 340 => b"00000_0000_01_000000000000", -- load, gr0
 341 => b"00000_0000_00_000000000001", -- 1
 342 => b"00001_0000_10_001000100111", -- store, gr0, P1BOMBACTIVE
 343 => b"00001_0011_10_001000100101", -- store, gr3, P1BOMBPOS
 344 => b"00000_0000_01_000000000000", -- load, gr0
 345 => b"00000_0000_00_000000010000", -- 16
 346 => b"00001_0000_10_001000100110", -- store, gr0, P1BOMBTIME
 347 => b"00000_0000_00_001000110001", -- load, gr0, BOMBS1
 348 => b"00010_0000_01_000000000000", -- add, gr0
 349 => b"00000_0000_00_000000000001", -- 1
 350 => b"00001_0000_10_001000110001", -- store, gr0, BOMBS1
 351 => b"00100_0000_01_000000000000", -- jump
 352 => b"00000_0000_00_000100111000", -- BTN1_R
 353 => b"00000_0000_00_001000110010", -- load, gr0, BOMBS2
 354 => b"00011_0000_00_001000110011", -- sub, gr0, MAXBOMBS
 355 => b"00110_0000_01_000000000000", -- beq
 356 => b"00000_0000_00_000100111010", -- BTN2_R
 357 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 358 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 359 => b"00000_0000_00_001000110111", -- load, gr0, YPOS2
 360 => b"01000_0000_01_000000000000", -- mul, gr0
 361 => b"00000_0000_00_000000001111", -- 15
 362 => b"00010_0000_00_001000110110", -- add, gr0, XPOS2
 363 => b"10000_0000_00_000000000000", -- tpoint, gr0
 364 => b"01111_0001_00_000000000000", -- tread, gr1
 365 => b"00011_0001_00_001000111111", -- sub, gr1, EGG
 366 => b"00110_0000_01_000000000000", -- beq
 367 => b"00000_0000_00_000100111010", -- BTN2_R
 368 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 369 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 370 => b"00000_0011_00_001000110111", -- load, gr3, YPOS2
 371 => b"00000_0010_00_001000111111", -- load, gr2, EGG
 372 => b"01000_0011_01_000000000000", -- mul, gr3
 373 => b"00000_0000_00_000000001111", -- 15
 374 => b"00010_0011_00_001000110110", -- add, gr3, XPOS2
 375 => b"10000_0011_00_000000000000", -- tpoint, gr3
 376 => b"01110_0010_00_000000000000", -- twrite, gr2
 377 => b"00000_0000_01_000000000000", -- load, gr0
 378 => b"00000_0000_00_000000000001", -- 1
 379 => b"00001_0000_10_001000101101", -- store, gr0, P2BOMBACTIVE
 380 => b"00001_0011_10_001000101011", -- store, gr3, P2BOMBPOS
 381 => b"00000_0000_01_000000000000", -- load, gr0
 382 => b"00000_0000_00_000000010000", -- 16
 383 => b"00001_0000_10_001000101100", -- store, gr0, P2BOMBTIME
 384 => b"00000_0000_00_001000110010", -- load, gr0, BOMBS2
 385 => b"00010_0000_01_000000000000", -- add, gr0
 386 => b"00000_0000_00_000000000001", -- 1
 387 => b"00001_0000_10_001000110010", -- store, gr0, BOMBS2
 388 => b"00100_0000_01_000000000000", -- jump
 389 => b"00000_0000_00_000100111010", -- BTN2_R
 390 => b"00000_0000_00_000000000000", -- 0
 391 => b"00100_0000_01_000000000000", -- jump
 392 => b"00000_0000_00_001000100011", -- COUNT1
 393 => b"10001_0000_01_000000000000", -- joy1r
 394 => b"00000_0000_00_000110011011", -- P1R
 395 => b"10011_0000_01_000000000000", -- joy1l
 396 => b"00000_0000_00_000110111101", -- P1L
 397 => b"10010_0000_01_000000000000", -- joy1u
 398 => b"00000_0000_00_000110101100", -- P1U
 399 => b"10100_0000_01_000000000000", -- joy1d
 400 => b"00000_0000_00_000111001110", -- P1D
 401 => b"10110_0000_01_000000000000", -- joy2r
 402 => b"00000_0000_00_000111011111", -- P2R
 403 => b"11000_0000_01_000000000000", -- joy2l
 404 => b"00000_0000_00_001000000001", -- P2L
 405 => b"10111_0000_01_000000000000", -- joy2u
 406 => b"00000_0000_00_000111110000", -- P2U
 407 => b"11001_0000_01_000000000000", -- joy2d
 408 => b"00000_0000_00_001000010010", -- P2D
 409 => b"00100_0000_01_000000000000", -- jump
 410 => b"00000_0000_00_000000000100", -- CONTROL_R
 411 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 412 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 413 => b"00000_0000_00_001000110101", -- load, gr0, YPOS1
 414 => b"01000_0000_01_000000000000", -- mul, gr0
 415 => b"00000_0000_00_000000001111", -- 15
 416 => b"00010_0000_00_001000110100", -- add, gr0, XPOS1
 417 => b"00010_0000_01_000000000000", -- add, gr0
 418 => b"00000_0000_00_000000000001", -- 1
 419 => b"10000_0000_00_000000000000", -- tpoint, gr0
 420 => b"01111_0001_00_000000000000", -- tread, gr1
 421 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 422 => b"00111_0000_01_000000000000", -- bne
 423 => b"00000_0000_00_000110001101", -- J1
 424 => b"00010_1100_01_000000000000", -- add, gr12
 425 => b"00000_0000_00_000000000001", -- 1
 426 => b"00100_0000_01_000000000000", -- jump
 427 => b"00000_0000_00_000110001101", -- J1
 428 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 429 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 430 => b"00000_0000_00_001000110101", -- load, gr0, YPOS1
 431 => b"00011_0000_01_000000000000", -- sub, gr0
 432 => b"00000_0000_00_000000000001", -- 1
 433 => b"01000_0000_01_000000000000", -- mul, gr0
 434 => b"00000_0000_00_000000001111", -- 15
 435 => b"00010_0000_00_001000110100", -- add, gr0, XPOS1
 436 => b"10000_0000_00_000000000000", -- tpoint, gr0
 437 => b"01111_0001_00_000000000000", -- tread, gr1
 438 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 439 => b"00111_0000_01_000000000000", -- bne
 440 => b"00000_0000_00_000110010001", -- J2
 441 => b"00011_1101_01_000000000000", -- sub, gr13
 442 => b"00000_0000_00_000000000001", -- 1
 443 => b"00100_0000_01_000000000000", -- jump
 444 => b"00000_0000_00_000110010001", -- J2
 445 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 446 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 447 => b"00000_0000_00_001000110101", -- load, gr0, YPOS1
 448 => b"01000_0000_01_000000000000", -- mul, gr0
 449 => b"00000_0000_00_000000001111", -- 15
 450 => b"00010_0000_00_001000110100", -- add, gr0, XPOS1
 451 => b"00011_0000_01_000000000000", -- sub, gr0
 452 => b"00000_0000_00_000000000001", -- 1
 453 => b"10000_0000_00_000000000000", -- tpoint, gr0
 454 => b"01111_0001_00_000000000000", -- tread, gr1
 455 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 456 => b"00111_0000_01_000000000000", -- bne
 457 => b"00000_0000_00_000110001101", -- J1
 458 => b"00011_1100_01_000000000000", -- sub, gr12
 459 => b"00000_0000_00_000000000001", -- 1
 460 => b"00100_0000_01_000000000000", -- jump
 461 => b"00000_0000_00_000110001101", -- J1
 462 => b"00001_1100_10_001000110100", -- store, gr12, XPOS1
 463 => b"00001_1101_10_001000110101", -- store, gr13, YPOS1
 464 => b"00000_0000_00_001000110101", -- load, gr0, YPOS1
 465 => b"00010_0000_01_000000000000", -- add, gr0
 466 => b"00000_0000_00_000000000001", -- 1
 467 => b"01000_0000_01_000000000000", -- mul, gr0
 468 => b"00000_0000_00_000000001111", -- 15
 469 => b"00010_0000_00_001000110100", -- add, gr0, XPOS1
 470 => b"10000_0000_00_000000000000", -- tpoint, gr0
 471 => b"01111_0001_00_000000000000", -- tread, gr1
 472 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 473 => b"00111_0000_01_000000000000", -- bne
 474 => b"00000_0000_00_000110010001", -- J2
 475 => b"00010_1101_01_000000000000", -- add, gr13
 476 => b"00000_0000_00_000000000001", -- 1
 477 => b"00100_0000_01_000000000000", -- jump
 478 => b"00000_0000_00_000110010001", -- J2
 479 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 480 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 481 => b"00000_0000_00_001000110111", -- load, gr0, YPOS2
 482 => b"01000_0000_01_000000000000", -- mul, gr0
 483 => b"00000_0000_00_000000001111", -- 15
 484 => b"00010_0000_00_001000110110", -- add, gr0, XPOS2
 485 => b"00010_0000_01_000000000000", -- add, gr0
 486 => b"00000_0000_00_000000000001", -- 1
 487 => b"10000_0000_00_000000000000", -- tpoint, gr0
 488 => b"01111_0001_00_000000000000", -- tread, gr1
 489 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 490 => b"00111_0000_01_000000000000", -- bne
 491 => b"00000_0000_00_000110010101", -- J3
 492 => b"00010_1110_01_000000000000", -- add, gr14
 493 => b"00000_0000_00_000000000001", -- 1
 494 => b"00100_0000_01_000000000000", -- jump
 495 => b"00000_0000_00_000110010101", -- J3
 496 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 497 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 498 => b"00000_0000_00_001000110111", -- load, gr0, YPOS2
 499 => b"00011_0000_01_000000000000", -- sub, gr0
 500 => b"00000_0000_00_000000000001", -- 1
 501 => b"01000_0000_01_000000000000", -- mul, gr0
 502 => b"00000_0000_00_000000001111", -- 15
 503 => b"00010_0000_00_001000110110", -- add, gr0, XPOS2
 504 => b"10000_0000_00_000000000000", -- tpoint, gr0
 505 => b"01111_0001_00_000000000000", -- tread, gr1
 506 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 507 => b"00111_0000_01_000000000000", -- bne
 508 => b"00000_0000_00_000000000100", -- CONTROL_R
 509 => b"00011_1111_01_000000000000", -- sub, gr15
 510 => b"00000_0000_00_000000000001", -- 1
 511 => b"00100_0000_01_000000000000", -- jump
 512 => b"00000_0000_00_000000000100", -- CONTROL_R
 513 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 514 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 515 => b"00000_0000_00_001000110111", -- load, gr0, YPOS2
 516 => b"01000_0000_01_000000000000", -- mul, gr0
 517 => b"00000_0000_00_000000001111", -- 15
 518 => b"00010_0000_00_001000110110", -- add, gr0, XPOS2
 519 => b"00011_0000_01_000000000000", -- sub, gr0
 520 => b"00000_0000_00_000000000001", -- 1
 521 => b"10000_0000_00_000000000000", -- tpoint, gr0
 522 => b"01111_0001_00_000000000000", -- tread, gr1
 523 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 524 => b"00111_0000_01_000000000000", -- bne
 525 => b"00000_0000_00_000110010101", -- J3
 526 => b"00011_1110_01_000000000000", -- sub, gr14
 527 => b"00000_0000_00_000000000001", -- 1
 528 => b"00100_0000_01_000000000000", -- jump
 529 => b"00000_0000_00_000110010101", -- J3
 530 => b"00001_1110_10_001000110110", -- store, gr14, XPOS2
 531 => b"00001_1111_10_001000110111", -- store, gr15, YPOS2
 532 => b"00000_0000_00_001000110111", -- load, gr0, YPOS2
 533 => b"00010_0000_01_000000000000", -- add, gr0
 534 => b"00000_0000_00_000000000001", -- 1
 535 => b"01000_0000_01_000000000000", -- mul, gr0
 536 => b"00000_0000_00_000000001111", -- 15
 537 => b"00010_0000_00_001000110110", -- add, gr0, XPOS2
 538 => b"10000_0000_00_000000000000", -- tpoint, gr0
 539 => b"01111_0001_00_000000000000", -- tread, gr1
 540 => b"00011_0001_00_001000111011", -- sub, gr1, GRASS
 541 => b"00111_0000_01_000000000000", -- bne
 542 => b"00000_0000_00_000000000100", -- CONTROL_R
 543 => b"00010_1111_01_000000000000", -- add, gr15
 544 => b"00000_0000_00_000000000001", -- 1
 545 => b"00100_0000_01_000000000000", -- jump
 546 => b"00000_0000_00_000000000100", -- CONTROL_R
 547 => b"00100_0000_01_000000000000", -- jump
 548 => b"00000_0000_00_000110001001", -- COUNT_R
 549 => b"00000_0000_00_000000000000", -- 0
 550 => b"00000_0000_00_000000000000", -- 0
 551 => b"00000_0000_00_000000000000", -- 0
 552 => b"00000_0000_00_000000000000", -- 0
 553 => b"00000_0000_00_000000000000", -- 0
 554 => b"00000_0000_00_000000000000", -- 0
 555 => b"00000_0000_00_000000000000", -- 0
 556 => b"00000_0000_00_000000000000", -- 0
 557 => b"00000_0000_00_000000000000", -- 0
 558 => b"00000_0000_00_000000000000", -- 0
 559 => b"00000_0000_00_000000000000", -- 0
 560 => b"00000_0000_00_000000000000", -- 0
 561 => b"00000_0000_00_000000000000", -- 0
 562 => b"00000_0000_00_000000000000", -- 0
 563 => b"00000_0000_00_000000000001", -- 1
 564 => b"00000_0000_00_000000000000", -- 0
 565 => b"00000_0000_00_000000000000", -- 0
 566 => b"00000_0000_00_000000000000", -- 0
 567 => b"00000_0000_00_000000000000", -- 0
 568 => b"00000_0000_00_000000000000", -- 0
 569 => b"00000_0000_00_000000000000", -- 0
 570 => b"00000_0000_00_000000000000", -- 0
 571 => b"00000_0000_00_000000000000", -- 0
 572 => b"00000_0000_00_000000000001", -- 1
 573 => b"00000_0000_00_000000000010", -- 2
 574 => b"00000_0000_00_000000000011", -- 3
 575 => b"00000_0000_00_000000000100", -- 4


    others => (others => 0)
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = 1 then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = 1 else PM(to_integer(pAddr));

end Behavioral; 
