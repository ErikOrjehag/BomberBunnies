library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

     0 => b"00000_1100_01_000000000000", -- load, gr12
   1 => b"00000_0000_00_000000000001", -- 1
   2 => b"00000_1110_01_000000000000", -- load, gr14
   3 => b"00000_0000_00_000000001101", -- 13
   4 => b"00000_1111_01_000000000000", -- load, gr15
   5 => b"00000_0000_00_000000001011", -- 11
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001110", -- EXPLOSION
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000010100010", -- CONTROL
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000001010111", -- BUTTON
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000000000110", -- MAIN
  14 => b"00000_0000_00_000100111101", -- load, gr0, MAIN_TIMER
  15 => b"00011_0000_01_000000000000", -- sub, gr0
  16 => b"00000_0000_00_000000101000", -- 40
  17 => b"00110_0000_01_000000000000", -- beq
  18 => b"00000_0000_00_000000011001", -- MAIN_TIMER_RESET
  19 => b"00000_0000_00_000100111101", -- load, gr0, MAIN_TIMER
  20 => b"00010_0000_01_000000000000", -- add, gr0
  21 => b"00000_0000_00_000000000001", -- 1
  22 => b"00001_0000_10_000100111101", -- store, gr0, MAIN_TIMER
  23 => b"00100_0000_01_000000000000", -- jump
  24 => b"00000_0000_00_000000001000", -- EXPLOSION_R
  25 => b"00000_0000_01_000000000000", -- load, gr0
  26 => b"00000_0000_00_000000000000", -- 0
  27 => b"00001_0000_10_000100111101", -- store, gr0, MAIN_TIMER
  28 => b"00000_0010_00_000100111110", -- load, gr2, BOMB11
  29 => b"00011_0010_01_000000000000", -- sub, gr2
  30 => b"00000_0000_00_000000000001", -- 1
  31 => b"00110_0000_01_000000000000", -- beq
  32 => b"00000_0000_00_000000001000", -- EXPLOSION_R
  33 => b"00000_0000_00_000101000100", -- load, gr0, TIMER11
  34 => b"00011_0000_01_000000000000", -- sub, gr0
  35 => b"00000_0000_00_111111111111", -- 4095
  36 => b"00110_0000_01_000000000000", -- beq
  37 => b"00000_0000_00_000000101010", -- BOMB11_EXPLOSION
  38 => b"00000_0000_00_000101000100", -- load, gr0, TIMER11
  39 => b"00010_0000_01_000000000000", -- add, gr0
  40 => b"00000_0000_00_000000000001", -- 1
  41 => b"00001_0000_10_000101000100", -- store, gr0, TIMER11
  42 => b"00000_0010_00_000101001010", -- load, gr2, BOMB11POS
  43 => b"00000_0011_00_000101010010", -- load, gr3, BOOM
  44 => b"10000_0010_00_000000000000", -- tpoint, gr2
  45 => b"01110_0011_00_000000000000", -- twrite, gr3
  46 => b"00010_0010_01_000000000000", -- add, gr2
  47 => b"00000_0000_00_000000000001", -- 1
  48 => b"10000_0010_00_000000000000", -- tpoint, gr2
  49 => b"01110_0011_00_000000000000", -- twrite, gr3
  50 => b"00010_0010_01_000000000000", -- add, gr2
  51 => b"00000_0000_00_000000000001", -- 1
  52 => b"10000_0010_00_000000000000", -- tpoint, gr2
  53 => b"01110_0011_00_000000000000", -- twrite, gr3
  54 => b"00000_0010_00_000101001010", -- load, gr2, BOMB11POS
  55 => b"00011_0010_01_000000000000", -- sub, gr2
  56 => b"00000_0000_00_000000000001", -- 1
  57 => b"10000_0010_00_000000000000", -- tpoint, gr2
  58 => b"01110_0011_00_000000000000", -- twrite, gr3
  59 => b"00011_0010_01_000000000000", -- sub, gr2
  60 => b"00000_0000_00_000000000001", -- 1
  61 => b"10000_0010_00_000000000000", -- tpoint, gr2
  62 => b"01110_0011_00_000000000000", -- twrite, gr3
  63 => b"00000_0010_00_000101001010", -- load, gr2, BOMB11POS
  64 => b"00010_0010_01_000000000000", -- add, gr2
  65 => b"00000_0000_00_000000001111", -- 15
  66 => b"10000_0010_00_000000000000", -- tpoint, gr2
  67 => b"01110_0011_00_000000000000", -- twrite, gr3
  68 => b"00010_0010_01_000000000000", -- add, gr2
  69 => b"00000_0000_00_000000001111", -- 15
  70 => b"10000_0010_00_000000000000", -- tpoint, gr2
  71 => b"01110_0011_00_000000000000", -- twrite, gr3
  72 => b"00000_0010_00_000101001010", -- load, gr2, BOMB11POS
  73 => b"00011_0010_01_000000000000", -- sub, gr2
  74 => b"00000_0000_00_000000001111", -- 15
  75 => b"10000_0010_00_000000000000", -- tpoint, gr2
  76 => b"01110_0011_00_000000000000", -- twrite, gr3
  77 => b"00011_0010_01_000000000000", -- sub, gr2
  78 => b"00000_0000_00_000000001111", -- 15
  79 => b"10000_0010_00_000000000000", -- tpoint, gr2
  80 => b"01110_0011_00_000000000000", -- twrite, gr3
  81 => b"00000_0000_01_000000000000", -- load, gr0
  82 => b"00000_0000_00_000000000000", -- 0
  83 => b"00001_0000_10_000100111110", -- store, gr0, BOMB11
  84 => b"00001_0000_10_000101000100", -- store, gr0, TIMER11
  85 => b"00100_0000_01_000000000000", -- jump
  86 => b"00000_0000_00_000000001000", -- EXPLOSION_R
  87 => b"10101_0000_01_000000000000", -- btn1
  88 => b"00000_0000_00_000001011101", -- BTN1
  89 => b"11010_0000_01_000000000000", -- btn2
  90 => b"00000_0000_00_000010000100", -- BTN2
  91 => b"00100_0000_01_000000000000", -- jump
  92 => b"00000_0000_00_000000001100", -- BUTTON_R
  93 => b"00000_0000_00_000101001100", -- load, gr0, BOMBCOUNT1
  94 => b"00011_0000_00_000101001110", -- sub, gr0, MAXBOMBS
  95 => b"00110_0000_01_000000000000", -- beq
  96 => b"00000_0000_00_000001011001", -- BTN1_R
  97 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
  98 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
  99 => b"00000_0000_00_000101010101", -- load, gr0, YPOS1
 100 => b"01000_0000_01_000000000000", -- mul, gr0
 101 => b"00000_0000_00_000000001111", -- 15
 102 => b"00010_0000_00_000101010100", -- add, gr0, XPOS1
 103 => b"10000_0000_00_000000000000", -- tpoint, gr0
 104 => b"01111_0001_00_000000000000", -- tread, gr1
 105 => b"00011_0001_00_000101010011", -- sub, gr1, EGG
 106 => b"00110_0000_01_000000000000", -- beq
 107 => b"00000_0000_00_000001011011", -- BTN2_R
 108 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
 109 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
 110 => b"00000_0011_00_000101010101", -- load, gr3, YPOS1
 111 => b"00000_0010_00_000101010011", -- load, gr2, EGG
 112 => b"01000_0011_01_000000000000", -- mul, gr3
 113 => b"00000_0000_00_000000001111", -- 15
 114 => b"00010_0011_00_000101010100", -- add, gr3, XPOS1
 115 => b"10000_0011_00_000000000000", -- tpoint, gr3
 116 => b"01110_0010_00_000000000000", -- twrite, gr2
 117 => b"00001_0011_10_000101001010", -- store, gr3, BOMB11POS
 118 => b"00000_0000_00_000101001100", -- load, gr0, BOMBCOUNT1
 119 => b"00010_0000_01_000000000000", -- add, gr0
 120 => b"00000_0000_00_000000000001", -- 1
 121 => b"00001_0000_10_000101001100", -- store, gr0, BOMBCOUNT1
 122 => b"00000_0000_00_000100111110", -- load, gr0, BOMB11
 123 => b"00011_0000_01_000000000000", -- sub, gr0
 124 => b"00000_0000_00_000000000001", -- 1
 125 => b"00110_0000_01_000000000000", -- beq
 126 => b"00000_0000_00_000001011001", -- BTN1_R
 127 => b"00010_0000_01_000000000000", -- add, gr0
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"00001_0000_10_000100111110", -- store, gr0, BOMB11
 130 => b"00100_0000_01_000000000000", -- jump
 131 => b"00000_0000_00_000001011001", -- BTN1_R
 132 => b"00000_0000_00_000101001101", -- load, gr0, BOMBCOUNT2
 133 => b"00011_0000_00_000101001110", -- sub, gr0, MAXBOMBS
 134 => b"00110_0000_01_000000000000", -- beq
 135 => b"00000_0000_00_000001011011", -- BTN2_R
 136 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 137 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 138 => b"00000_0000_00_000101010111", -- load, gr0, YPOS2
 139 => b"01000_0000_01_000000000000", -- mul, gr0
 140 => b"00000_0000_00_000000001111", -- 15
 141 => b"00010_0000_00_000101010110", -- add, gr0, XPOS2
 142 => b"10000_0000_00_000000000000", -- tpoint, gr0
 143 => b"01111_0001_00_000000000000", -- tread, gr1
 144 => b"00011_0001_00_000101010011", -- sub, gr1, EGG
 145 => b"00110_0000_01_000000000000", -- beq
 146 => b"00000_0000_00_000001011011", -- BTN2_R
 147 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 148 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 149 => b"00000_0011_00_000101010111", -- load, gr3, YPOS2
 150 => b"00000_0010_00_000101010011", -- load, gr2, EGG
 151 => b"01000_0011_01_000000000000", -- mul, gr3
 152 => b"00000_0000_00_000000001111", -- 15
 153 => b"00010_0011_00_000101010110", -- add, gr3, XPOS2
 154 => b"10000_0011_00_000000000000", -- tpoint, gr3
 155 => b"01110_0010_00_000000000000", -- twrite, gr2
 156 => b"00000_0000_00_000101001101", -- load, gr0, BOMBCOUNT2
 157 => b"00010_0000_01_000000000000", -- add, gr0
 158 => b"00000_0000_00_000000000001", -- 1
 159 => b"00001_0000_10_000101001101", -- store, gr0, BOMBCOUNT2
 160 => b"00100_0000_01_000000000000", -- jump
 161 => b"00000_0000_00_000001011011", -- BTN2_R
 162 => b"10001_0000_01_000000000000", -- joy1r
 163 => b"00000_0000_00_000010110100", -- P1R
 164 => b"10011_0000_01_000000000000", -- joy1l
 165 => b"00000_0000_00_000011010110", -- P1L
 166 => b"10010_0000_01_000000000000", -- joy1u
 167 => b"00000_0000_00_000011000101", -- P1U
 168 => b"10100_0000_01_000000000000", -- joy1d
 169 => b"00000_0000_00_000011100111", -- P1D
 170 => b"10110_0000_01_000000000000", -- joy2r
 171 => b"00000_0000_00_000011111000", -- P2R
 172 => b"11000_0000_01_000000000000", -- joy2l
 173 => b"00000_0000_00_000100011010", -- P2L
 174 => b"10111_0000_01_000000000000", -- joy2u
 175 => b"00000_0000_00_000100001001", -- P2U
 176 => b"11001_0000_01_000000000000", -- joy2d
 177 => b"00000_0000_00_000100101011", -- P2D
 178 => b"00100_0000_01_000000000000", -- jump
 179 => b"00000_0000_00_000000001010", -- CONTROL_R
 180 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
 181 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
 182 => b"00000_0000_00_000101010101", -- load, gr0, YPOS1
 183 => b"01000_0000_01_000000000000", -- mul, gr0
 184 => b"00000_0000_00_000000001111", -- 15
 185 => b"00010_0000_00_000101010100", -- add, gr0, XPOS1
 186 => b"00010_0000_01_000000000000", -- add, gr0
 187 => b"00000_0000_00_000000000001", -- 1
 188 => b"10000_0000_00_000000000000", -- tpoint, gr0
 189 => b"01111_0001_00_000000000000", -- tread, gr1
 190 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000010100110", -- J1
 193 => b"00010_1100_01_000000000000", -- add, gr12
 194 => b"00000_0000_00_000000000001", -- 1
 195 => b"00100_0000_01_000000000000", -- jump
 196 => b"00000_0000_00_000010100110", -- J1
 197 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
 198 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
 199 => b"00000_0000_00_000101010101", -- load, gr0, YPOS1
 200 => b"00011_0000_01_000000000000", -- sub, gr0
 201 => b"00000_0000_00_000000000001", -- 1
 202 => b"01000_0000_01_000000000000", -- mul, gr0
 203 => b"00000_0000_00_000000001111", -- 15
 204 => b"00010_0000_00_000101010100", -- add, gr0, XPOS1
 205 => b"10000_0000_00_000000000000", -- tpoint, gr0
 206 => b"01111_0001_00_000000000000", -- tread, gr1
 207 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 208 => b"00111_0000_01_000000000000", -- bne
 209 => b"00000_0000_00_000010101010", -- J2
 210 => b"00011_1101_01_000000000000", -- sub, gr13
 211 => b"00000_0000_00_000000000001", -- 1
 212 => b"00100_0000_01_000000000000", -- jump
 213 => b"00000_0000_00_000010101010", -- J2
 214 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
 215 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
 216 => b"00000_0000_00_000101010101", -- load, gr0, YPOS1
 217 => b"01000_0000_01_000000000000", -- mul, gr0
 218 => b"00000_0000_00_000000001111", -- 15
 219 => b"00010_0000_00_000101010100", -- add, gr0, XPOS1
 220 => b"00011_0000_01_000000000000", -- sub, gr0
 221 => b"00000_0000_00_000000000001", -- 1
 222 => b"10000_0000_00_000000000000", -- tpoint, gr0
 223 => b"01111_0001_00_000000000000", -- tread, gr1
 224 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 225 => b"00111_0000_01_000000000000", -- bne
 226 => b"00000_0000_00_000010100110", -- J1
 227 => b"00011_1100_01_000000000000", -- sub, gr12
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00100_0000_01_000000000000", -- jump
 230 => b"00000_0000_00_000010100110", -- J1
 231 => b"00001_1100_10_000101010100", -- store, gr12, XPOS1
 232 => b"00001_1101_10_000101010101", -- store, gr13, YPOS1
 233 => b"00000_0000_00_000101010101", -- load, gr0, YPOS1
 234 => b"00010_0000_01_000000000000", -- add, gr0
 235 => b"00000_0000_00_000000000001", -- 1
 236 => b"01000_0000_01_000000000000", -- mul, gr0
 237 => b"00000_0000_00_000000001111", -- 15
 238 => b"00010_0000_00_000101010100", -- add, gr0, XPOS1
 239 => b"10000_0000_00_000000000000", -- tpoint, gr0
 240 => b"01111_0001_00_000000000000", -- tread, gr1
 241 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 242 => b"00111_0000_01_000000000000", -- bne
 243 => b"00000_0000_00_000010101010", -- J2
 244 => b"00010_1101_01_000000000000", -- add, gr13
 245 => b"00000_0000_00_000000000001", -- 1
 246 => b"00100_0000_01_000000000000", -- jump
 247 => b"00000_0000_00_000010101010", -- J2
 248 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 249 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 250 => b"00000_0000_00_000101010111", -- load, gr0, YPOS2
 251 => b"01000_0000_01_000000000000", -- mul, gr0
 252 => b"00000_0000_00_000000001111", -- 15
 253 => b"00010_0000_00_000101010110", -- add, gr0, XPOS2
 254 => b"00010_0000_01_000000000000", -- add, gr0
 255 => b"00000_0000_00_000000000001", -- 1
 256 => b"10000_0000_00_000000000000", -- tpoint, gr0
 257 => b"01111_0001_00_000000000000", -- tread, gr1
 258 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 259 => b"00111_0000_01_000000000000", -- bne
 260 => b"00000_0000_00_000010101110", -- J3
 261 => b"00010_1110_01_000000000000", -- add, gr14
 262 => b"00000_0000_00_000000000001", -- 1
 263 => b"00100_0000_01_000000000000", -- jump
 264 => b"00000_0000_00_000010101110", -- J3
 265 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 266 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 267 => b"00000_0000_00_000101010111", -- load, gr0, YPOS2
 268 => b"00011_0000_01_000000000000", -- sub, gr0
 269 => b"00000_0000_00_000000000001", -- 1
 270 => b"01000_0000_01_000000000000", -- mul, gr0
 271 => b"00000_0000_00_000000001111", -- 15
 272 => b"00010_0000_00_000101010110", -- add, gr0, XPOS2
 273 => b"10000_0000_00_000000000000", -- tpoint, gr0
 274 => b"01111_0001_00_000000000000", -- tread, gr1
 275 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 276 => b"00111_0000_01_000000000000", -- bne
 277 => b"00000_0000_00_000000001010", -- CONTROL_R
 278 => b"00011_1111_01_000000000000", -- sub, gr15
 279 => b"00000_0000_00_000000000001", -- 1
 280 => b"00100_0000_01_000000000000", -- jump
 281 => b"00000_0000_00_000000001010", -- CONTROL_R
 282 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 283 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 284 => b"00000_0000_00_000101010111", -- load, gr0, YPOS2
 285 => b"01000_0000_01_000000000000", -- mul, gr0
 286 => b"00000_0000_00_000000001111", -- 15
 287 => b"00010_0000_00_000101010110", -- add, gr0, XPOS2
 288 => b"00011_0000_01_000000000000", -- sub, gr0
 289 => b"00000_0000_00_000000000001", -- 1
 290 => b"10000_0000_00_000000000000", -- tpoint, gr0
 291 => b"01111_0001_00_000000000000", -- tread, gr1
 292 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 293 => b"00111_0000_01_000000000000", -- bne
 294 => b"00000_0000_00_000010101110", -- J3
 295 => b"00011_1110_01_000000000000", -- sub, gr14
 296 => b"00000_0000_00_000000000001", -- 1
 297 => b"00100_0000_01_000000000000", -- jump
 298 => b"00000_0000_00_000010101110", -- J3
 299 => b"00001_1110_10_000101010110", -- store, gr14, XPOS2
 300 => b"00001_1111_10_000101010111", -- store, gr15, YPOS2
 301 => b"00000_0000_00_000101010111", -- load, gr0, YPOS2
 302 => b"00010_0000_01_000000000000", -- add, gr0
 303 => b"00000_0000_00_000000000001", -- 1
 304 => b"01000_0000_01_000000000000", -- mul, gr0
 305 => b"00000_0000_00_000000001111", -- 15
 306 => b"00010_0000_00_000101010110", -- add, gr0, XPOS2
 307 => b"10000_0000_00_000000000000", -- tpoint, gr0
 308 => b"01111_0001_00_000000000000", -- tread, gr1
 309 => b"00011_0001_00_000101001111", -- sub, gr1, GRASS
 310 => b"00111_0000_01_000000000000", -- bne
 311 => b"00000_0000_00_000000001010", -- CONTROL_R
 312 => b"00010_1111_01_000000000000", -- add, gr15
 313 => b"00000_0000_00_000000000001", -- 1
 314 => b"00100_0000_01_000000000000", -- jump
 315 => b"00000_0000_00_000000001010", -- CONTROL_R
 316 => b"00000_0000_00_000000000000", -- 0
 317 => b"00000_0000_00_000000000000", -- 0
 318 => b"00000_0000_00_000000000000", -- 0
 319 => b"00000_0000_00_000000000000", -- 0
 320 => b"00000_0000_00_000000000000", -- 0
 321 => b"00000_0000_00_000000000000", -- 0
 322 => b"00000_0000_00_000000000000", -- 0
 323 => b"00000_0000_00_000000000000", -- 0
 324 => b"00000_0000_00_000000000000", -- 0
 325 => b"00000_0000_00_000000000000", -- 0
 326 => b"00000_0000_00_000000000000", -- 0
 327 => b"00000_0000_00_000000000000", -- 0
 328 => b"00000_0000_00_000000000000", -- 0
 329 => b"00000_0000_00_000000000000", -- 0
 330 => b"00000_0000_00_000000000000", -- 0
 331 => b"00000_0000_00_000000000000", -- 0
 332 => b"00000_0000_00_000000000000", -- 0
 333 => b"00000_0000_00_000000000000", -- 0
 334 => b"00000_0000_00_000000000011", -- 3
 335 => b"00000_0000_00_000000000000", -- 0
 336 => b"00000_0000_00_000000000001", -- 1
 337 => b"00000_0000_00_000000000010", -- 2
 338 => b"00000_0000_00_000000000011", -- 3
 339 => b"00000_0000_00_000000000100", -- 4
 340 => b"00000_0000_00_000000000000", -- 0
 341 => b"00000_0000_00_000000000000", -- 0
 342 => b"00000_0000_00_000000000000", -- 0
 343 => b"00000_0000_00_000000000000", -- 0



    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral;


