library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity MICRO_MEMORY is
  port (
    uAddr : in unsigned(8 downto 0);
    uData : out std_logic_vector(29 downto 0));
end MICRO_MEMORY;

architecture Behavioral of MICRO_MEMORY is

-- micro Memory
type u_mem_t is array (0 to 511) of std_logic_vector(29 downto 0);
constant u_mem_c : u_mem_t := (
  -- AR 0110
       --  ALU   TB   FB  S P LC  SEQ  uADR
    0 => b"0000_0100_0001_0_0_00_0000_000000000",  -- H�mtfas
    1 => b"0000_0011_0010_0_1_00_0000_000000000",
    
    2 => b"0000_0000_0000_0_0_00_0010_000000000",  -- Start
    
    3 => b"0000_0010_0001_0_0_00_0001_000000000",  -- Direktadressering
    
    4 => b"0000_0100_0001_0_1_00_0001_000000000",  -- Immediate
    
    5 => b"0000_0010_0001_0_0_00_0000_000000000",  -- Indirekt adressering
    6 => b"0000_0011_0001_0_0_00_0001_000000000",
    
    7 => b"0000_0110_0000_0_0_00_0000_000000000",  -- Indexerad adressering
    8 => b"1000_0101_0000_0_0_00_0000_000000000",
    9 => b"0000_0110_0001_0_0_00_0001_000000000",
    
    
    10 => b"0000_0011_0101_0_0_00_0011_000000000",  -- LOAD (GRx, M, ADDR)
    
    11 => b"0000_0101_0011_0_0_00_0011_000000000",  -- STORE (GRx, M, ADDR)
    
    12 => b"0001_0011_0000_0_0_00_0000_000000000",  -- ADD (GRx, M, ADDR)
    13 => b"0100_0101_0000_0_0_00_0000_000000000",
    14 => b"0000_0110_0101_0_0_00_0011_000000000",
    
    15 => b"0001_0101_0000_0_0_00_0000_000000000",  -- SUB (GRx, M, ADDR)
    16 => b"0101_0011_0000_0_0_00_0000_000000000",
    17 => b"0000_0110_0101_0_0_00_0011_000000000",
    
    18 => b"0000_0011_0100_0_0_00_0011_000000000",  -- JUMP
    
    19 => b"0000_0011_0000_0_0_00_0000_000000000",  -- SLEEP
    20 => b"0000_0000_0000_0_0_10_0000_000000000",
    21 => b"0000_0000_0000_0_0_01_0000_000000000",
    22 => b"0000_0000_0000_0_0_00_1100_000010101",
    23 => b"0000_0000_0000_0_0_00_0011_000000000",

    24 => b"0000_0000_0000_0_0_00_1000_000010010",  -- BEQ (g�r till JUMP om z=1)
    25 => b"0000_0000_0000_0_0_00_0011_000000000",

    26 => b"0000_0000_0000_0_0_00_0100_000010010",  -- BNE (g�r till JUMP om z=0 annars PC+1)
    27 => b"0000_0000_0000_0_1_00_0011_000000000",

    28 => b"0000_1010_0101_0_0_00_0011_000000000",  -- JOY1X

    29 => b"0000_1011_0101_0_0_00_0011_000000000",  -- JOY1Y

    30 => b"0000_1100_0101_0_0_00_0011_000000000",  -- BTN1

    31 => b"0000_1101_0101_0_0_00_0011_000000000",  -- JOY2X

    32 => b"0000_1110_0101_0_0_00_0011_000000000",  -- JOY2Y

    33 => b"0000_1111_0101_0_0_00_0011_000000000",  -- BTN2

    34 => b"0000_0101_1000_0_0_00_0101_000000000",  -- GRx till tileWrite,
    35 => b"0000_0000_0000_0_0_00_0011_000000000",

    36 => b"0000_1000_0101_0_0_00_0110_000000000",  -- tileRead to GRx
    37 => b"0000_0000_0000_0_0_00_0011_000000000",

    38 => b"0000_0101_1001_0_0_00_0011_000000000",  -- GRx to tilePointer
    
    others => (others => '0')
  );

signal uMem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= uMem(to_integer(uAddr));

end Behavioral;
