library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PROGRAM_MEMORY is
  
  port (
    clk : in std_logic;
    pAddr : in  unsigned(11 downto 0);
    PM_out : out std_logic_vector(22 downto 0);
    PM_in : in std_logic_vector(22 downto 0);
    PM_write : in std_logic
    );
  
end PROGRAM_MEMORY;

architecture Behavioral of PROGRAM_MEMORY is

  -- Add names for different operations that are binary?
  -- operations
  constant load : std_logic_vector        := "00000";
  constant store : std_logic_vector       := "00001";
  constant add : std_logic_vector         := "00010";
  constant sub : std_logic_vector         := "00011";
  constant jump : std_logic_vector        := "00100";
  constant sleep : std_logic_vector       := "00101";
  constant beq : std_logic_vector         := "00110";
  constant bne : std_logic_vector         := "00111";
  constant tileWrite : std_logic_vector   := "01110";
  constant tileRead : std_logic_vector    := "01111";
  constant tilePointer : std_logic_vector := "10000";
  constant joy1r : std_logic_vector       := "10001";
  constant joy1u : std_logic_vector       := "10010";
  constant joy1l : std_logic_vector       := "10011";
  constant joy1d : std_logic_vector       := "10100";
  constant btn1 : std_logic_vector        := "10101";
  constant joy2r : std_logic_vector       := "10110";
  constant joy2u : std_logic_vector       := "10111";
  constant joy2l : std_logic_vector       := "11000";
  constant joy2d : std_logic_vector       := "11001";
  constant btn2 : std_logic_vector        := "11010";

  -- GRx
  constant gr0 : std_logic_vector  := "0000";
  constant gr1 : std_logic_vector  := "0001";
  constant gr2 : std_logic_vector  := "0010";
  constant gr3 : std_logic_vector  := "0011";
  constant gr4 : std_logic_vector  := "0100";
  constant gr5 : std_logic_vector  := "0101";
  constant gr6 : std_logic_vector  := "0110";
  constant gr7 : std_logic_vector  := "0111";
  constant gr8 : std_logic_vector  := "1000";
  constant gr9 : std_logic_vector  := "1001";
  constant gr10 : std_logic_vector := "1010";
  constant gr11 : std_logic_vector := "1011";
  constant gr12 : std_logic_vector := "1100";
  constant gr13 : std_logic_vector := "1101";
  constant gr14 : std_logic_vector := "1110";
  constant gr15 : std_logic_vector := "1111";

  -- Program memory
  type pm_t is array (0 to 2047) of std_logic_vector(22 downto 0);  --2047
  constant pm_c : pm_t := (
       -- OP    GRx  M  Adr

   0 => b"00100_0000_01_000000000000", -- jump
   1 => b"00000_0000_00_001001001110", -- CONTROL
   2 => b"00100_0000_01_000000000000", -- jump
   3 => b"00000_0000_00_000110010100", -- BUTTON
   4 => b"00100_0000_01_000000000000", -- jump
   5 => b"00000_0000_00_000011000100", -- TICKBOMBS
   6 => b"00100_0000_01_000000000000", -- jump
   7 => b"00000_0000_00_000000001010", -- TICKEXPLOSIONS
   8 => b"00100_0000_01_000000000000", -- jump
   9 => b"00000_0000_00_000000000000", -- MAIN
  10 => b"00100_0000_01_000000000000", -- jump
  11 => b"00000_0000_00_000000010000", -- BOOM1
  12 => b"00100_0000_01_000000000000", -- jump
  13 => b"00000_0000_00_000001101010", -- BOOM2
  14 => b"00100_0000_01_000000000000", -- jump
  15 => b"00000_0000_00_000000001000", -- TICKEXPLOSIONS_R
  16 => b"00000_0000_00_001011110000", -- load, gr0, P1EXPLOSION1ACTIVE
  17 => b"00011_0000_01_000000000000", -- sub, gr0
  18 => b"00000_0000_00_000000000001", -- 1
  19 => b"00111_0000_01_000000000000", -- bne
  20 => b"00000_0000_00_000000001100", -- BOOM1_R
  21 => b"00000_0000_00_001011101111", -- load, gr0, P1EXPLOSION1TIME
  22 => b"00011_0000_01_000000000000", -- sub, gr0
  23 => b"00000_0000_00_000000000001", -- 1
  24 => b"00001_0000_10_001011101111", -- store, gr0, P1EXPLOSION1TIME
  25 => b"00000_0000_00_001011101111", -- load, gr0, P1EXPLOSION1TIME
  26 => b"00011_0000_01_000000000000", -- sub, gr0
  27 => b"00000_0000_00_000000000000", -- 0
  28 => b"00111_0000_01_000000000000", -- bne
  29 => b"00000_0000_00_000000001100", -- BOOM1_R
  30 => b"00000_0000_01_000000000000", -- load, gr0
  31 => b"00000_0000_00_000000000000", -- 0
  32 => b"00001_0000_10_001011110000", -- store, gr0, P1EXPLOSION1ACTIVE
  33 => b"00000_0010_00_001011110001", -- load, gr2, P1EXPLOSION1POS
  34 => b"00000_0011_00_001100011010", -- load, gr3, GRASS
  35 => b"10000_0010_00_000000000000", -- tpoint, gr2
  36 => b"01110_0011_00_000000000000", -- twrite, gr3
  37 => b"00010_0010_01_000000000000", -- add, gr2
  38 => b"00000_0000_00_000000000001", -- 1
  39 => b"10000_0010_00_000000000000", -- tpoint, gr2
  40 => b"01111_0000_00_000000000000", -- tread, gr0
  41 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  42 => b"00111_0000_01_000000000000", -- bne
  43 => b"00000_0000_00_000000110101", -- E1LEFT
  44 => b"01110_0011_00_000000000000", -- twrite, gr3
  45 => b"00010_0010_01_000000000000", -- add, gr2
  46 => b"00000_0000_00_000000000001", -- 1
  47 => b"10000_0010_00_000000000000", -- tpoint, gr2
  48 => b"01111_0000_00_000000000000", -- tread, gr0
  49 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  50 => b"00111_0000_01_000000000000", -- bne
  51 => b"00000_0000_00_000000110101", -- E1LEFT
  52 => b"01110_0011_00_000000000000", -- twrite, gr3
  53 => b"00000_0010_00_001011110001", -- load, gr2, P1EXPLOSION1POS
  54 => b"00011_0010_01_000000000000", -- sub, gr2
  55 => b"00000_0000_00_000000000001", -- 1
  56 => b"10000_0010_00_000000000000", -- tpoint, gr2
  57 => b"01111_0000_00_000000000000", -- tread, gr0
  58 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  59 => b"00111_0000_01_000000000000", -- bne
  60 => b"00000_0000_00_000001000110", -- E1DOWN
  61 => b"01110_0011_00_000000000000", -- twrite, gr3
  62 => b"00011_0010_01_000000000000", -- sub, gr2
  63 => b"00000_0000_00_000000000001", -- 1
  64 => b"10000_0010_00_000000000000", -- tpoint, gr2
  65 => b"01111_0000_00_000000000000", -- tread, gr0
  66 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  67 => b"00111_0000_01_000000000000", -- bne
  68 => b"00000_0000_00_000001000110", -- E1DOWN
  69 => b"01110_0011_00_000000000000", -- twrite, gr3
  70 => b"00000_0010_00_001011110001", -- load, gr2, P1EXPLOSION1POS
  71 => b"00010_0010_01_000000000000", -- add, gr2
  72 => b"00000_0000_00_000000001111", -- 15
  73 => b"10000_0010_00_000000000000", -- tpoint, gr2
  74 => b"01111_0000_00_000000000000", -- tread, gr0
  75 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  76 => b"00111_0000_01_000000000000", -- bne
  77 => b"00000_0000_00_000001010111", -- E1UP
  78 => b"01110_0011_00_000000000000", -- twrite, gr3
  79 => b"00010_0010_01_000000000000", -- add, gr2
  80 => b"00000_0000_00_000000001111", -- 15
  81 => b"10000_0010_00_000000000000", -- tpoint, gr2
  82 => b"01111_0000_00_000000000000", -- tread, gr0
  83 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  84 => b"00111_0000_01_000000000000", -- bne
  85 => b"00000_0000_00_000001010111", -- E1UP
  86 => b"01110_0011_00_000000000000", -- twrite, gr3
  87 => b"00000_0010_00_001011110001", -- load, gr2, P1EXPLOSION1POS
  88 => b"00011_0010_01_000000000000", -- sub, gr2
  89 => b"00000_0000_00_000000001111", -- 15
  90 => b"10000_0010_00_000000000000", -- tpoint, gr2
  91 => b"01111_0000_00_000000000000", -- tread, gr0
  92 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
  93 => b"00111_0000_01_000000000000", -- bne
  94 => b"00000_0000_00_000000001100", -- BOOM1_R
  95 => b"01110_0011_00_000000000000", -- twrite, gr3
  96 => b"00011_0010_01_000000000000", -- sub, gr2
  97 => b"00000_0000_00_000000001111", -- 15
  98 => b"10000_0010_00_000000000000", -- tpoint, gr2
  99 => b"01111_0000_00_000000000000", -- tread, gr0
 100 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 101 => b"00111_0000_01_000000000000", -- bne
 102 => b"00000_0000_00_000000001100", -- BOOM1_R
 103 => b"01110_0011_00_000000000000", -- twrite, gr3
 104 => b"00100_0000_01_000000000000", -- jump
 105 => b"00000_0000_00_000000001100", -- BOOM1_R
 106 => b"00000_0000_00_001100000010", -- load, gr0, P2EXPLOSION1ACTIVE
 107 => b"00011_0000_01_000000000000", -- sub, gr0
 108 => b"00000_0000_00_000000000001", -- 1
 109 => b"00111_0000_01_000000000000", -- bne
 110 => b"00000_0000_00_000000001110", -- BOOM2_R
 111 => b"00000_0000_00_001100000001", -- load, gr0, P2EXPLOSION1TIME
 112 => b"00011_0000_01_000000000000", -- sub, gr0
 113 => b"00000_0000_00_000000000001", -- 1
 114 => b"00001_0000_10_001100000001", -- store, gr0, P2EXPLOSION1TIME
 115 => b"00000_0000_00_001100000001", -- load, gr0, P2EXPLOSION1TIME
 116 => b"00011_0000_01_000000000000", -- sub, gr0
 117 => b"00000_0000_00_000000000000", -- 0
 118 => b"00111_0000_01_000000000000", -- bne
 119 => b"00000_0000_00_000000001110", -- BOOM2_R
 120 => b"00000_0000_01_000000000000", -- load, gr0
 121 => b"00000_0000_00_000000000000", -- 0
 122 => b"00001_0000_10_001100000010", -- store, gr0, P2EXPLOSION1ACTIVE
 123 => b"00000_0010_00_001100000011", -- load, gr2, P2EXPLOSION1POS
 124 => b"00000_0011_00_001100011010", -- load, gr3, GRASS
 125 => b"10000_0010_00_000000000000", -- tpoint, gr2
 126 => b"01110_0011_00_000000000000", -- twrite, gr3
 127 => b"00010_0010_01_000000000000", -- add, gr2
 128 => b"00000_0000_00_000000000001", -- 1
 129 => b"10000_0010_00_000000000000", -- tpoint, gr2
 130 => b"01111_0000_00_000000000000", -- tread, gr0
 131 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 132 => b"00111_0000_01_000000000000", -- bne
 133 => b"00000_0000_00_000010001111", -- E2LEFT
 134 => b"01110_0011_00_000000000000", -- twrite, gr3
 135 => b"00010_0010_01_000000000000", -- add, gr2
 136 => b"00000_0000_00_000000000001", -- 1
 137 => b"10000_0010_00_000000000000", -- tpoint, gr2
 138 => b"01111_0000_00_000000000000", -- tread, gr0
 139 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 140 => b"00111_0000_01_000000000000", -- bne
 141 => b"00000_0000_00_000010001111", -- E2LEFT
 142 => b"01110_0011_00_000000000000", -- twrite, gr3
 143 => b"00000_0010_00_001100000011", -- load, gr2, P2EXPLOSION1POS
 144 => b"00011_0010_01_000000000000", -- sub, gr2
 145 => b"00000_0000_00_000000000001", -- 1
 146 => b"10000_0010_00_000000000000", -- tpoint, gr2
 147 => b"01111_0000_00_000000000000", -- tread, gr0
 148 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 149 => b"00111_0000_01_000000000000", -- bne
 150 => b"00000_0000_00_000010100000", -- E2DOWN
 151 => b"01110_0011_00_000000000000", -- twrite, gr3
 152 => b"00011_0010_01_000000000000", -- sub, gr2
 153 => b"00000_0000_00_000000000001", -- 1
 154 => b"10000_0010_00_000000000000", -- tpoint, gr2
 155 => b"01111_0000_00_000000000000", -- tread, gr0
 156 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 157 => b"00111_0000_01_000000000000", -- bne
 158 => b"00000_0000_00_000010100000", -- E2DOWN
 159 => b"01110_0011_00_000000000000", -- twrite, gr3
 160 => b"00000_0010_00_001100000011", -- load, gr2, P2EXPLOSION1POS
 161 => b"00010_0010_01_000000000000", -- add, gr2
 162 => b"00000_0000_00_000000001111", -- 15
 163 => b"10000_0010_00_000000000000", -- tpoint, gr2
 164 => b"01111_0000_00_000000000000", -- tread, gr0
 165 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 166 => b"00111_0000_01_000000000000", -- bne
 167 => b"00000_0000_00_000010110001", -- E2UP
 168 => b"01110_0011_00_000000000000", -- twrite, gr3
 169 => b"00010_0010_01_000000000000", -- add, gr2
 170 => b"00000_0000_00_000000001111", -- 15
 171 => b"10000_0010_00_000000000000", -- tpoint, gr2
 172 => b"01111_0000_00_000000000000", -- tread, gr0
 173 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 174 => b"00111_0000_01_000000000000", -- bne
 175 => b"00000_0000_00_000010110001", -- E2UP
 176 => b"01110_0011_00_000000000000", -- twrite, gr3
 177 => b"00000_0010_00_001100000011", -- load, gr2, P2EXPLOSION1POS
 178 => b"00011_0010_01_000000000000", -- sub, gr2
 179 => b"00000_0000_00_000000001111", -- 15
 180 => b"10000_0010_00_000000000000", -- tpoint, gr2
 181 => b"01111_0000_00_000000000000", -- tread, gr0
 182 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 183 => b"00111_0000_01_000000000000", -- bne
 184 => b"00000_0000_00_000000001110", -- BOOM2_R
 185 => b"01110_0011_00_000000000000", -- twrite, gr3
 186 => b"00011_0010_01_000000000000", -- sub, gr2
 187 => b"00000_0000_00_000000001111", -- 15
 188 => b"10000_0010_00_000000000000", -- tpoint, gr2
 189 => b"01111_0000_00_000000000000", -- tread, gr0
 190 => b"00011_0000_00_001100011101", -- sub, gr0, EXPLOSION
 191 => b"00111_0000_01_000000000000", -- bne
 192 => b"00000_0000_00_000000001110", -- BOOM2_R
 193 => b"01110_0011_00_000000000000", -- twrite, gr3
 194 => b"00100_0000_01_000000000000", -- jump
 195 => b"00000_0000_00_000000001110", -- BOOM2_R
 196 => b"00100_0000_01_000000000000", -- jump
 197 => b"00000_0000_00_000011001010", -- TICKBOMB1
 198 => b"00100_0000_01_000000000000", -- jump
 199 => b"00000_0000_00_000100101111", -- TICKBOMB2
 200 => b"00100_0000_01_000000000000", -- jump
 201 => b"00000_0000_00_000000000110", -- TICKBOMBS_R
 202 => b"00000_0000_00_001011101110", -- load, gr0, P1BOMB1ACTIVE
 203 => b"00011_0000_01_000000000000", -- sub, gr0
 204 => b"00000_0000_00_000000000001", -- 1
 205 => b"00111_0000_01_000000000000", -- bne
 206 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 207 => b"00000_0000_00_001011101101", -- load, gr0, P1BOMB1TIME
 208 => b"00011_0000_01_000000000000", -- sub, gr0
 209 => b"00000_0000_00_000000000001", -- 1
 210 => b"00001_0000_10_001011101101", -- store, gr0, P1BOMB1TIME
 211 => b"00000_0000_01_000000000000", -- load, gr0
 212 => b"00000_0000_00_000000000000", -- 0
 213 => b"00011_0000_00_001011101101", -- sub, gr0, P1BOMB1TIME
 214 => b"00110_0000_01_000000000000", -- beq
 215 => b"00000_0000_00_000011011010", -- EXPLODE1
 216 => b"00100_0000_01_000000000000", -- jump
 217 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 218 => b"00000_0000_00_001011101100", -- load, gr0, P1BOMB1POS
 219 => b"00001_0000_10_001011110001", -- store, gr0, P1EXPLOSION1POS
 220 => b"00000_0000_01_000000000000", -- load, gr0
 221 => b"00000_0000_00_000000000001", -- 1
 222 => b"00001_0000_10_001011110000", -- store, gr0, P1EXPLOSION1ACTIVE
 223 => b"00000_0000_01_000000000000", -- load, gr0
 224 => b"00000_0000_00_000000000010", -- 2
 225 => b"00001_0000_10_001011101111", -- store, gr0, P1EXPLOSION1TIME
 226 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 227 => b"00011_0000_01_000000000000", -- sub, gr0
 228 => b"00000_0000_00_000000000001", -- 1
 229 => b"00001_0000_10_001100010000", -- store, gr0, P1BOMBCOUNT
 230 => b"00000_0010_00_001011101100", -- load, gr2, P1BOMB1POS
 231 => b"00000_0011_00_001100011101", -- load, gr3, EXPLOSION
 232 => b"10000_0010_00_000000000000", -- tpoint, gr2
 233 => b"01110_0011_00_000000000000", -- twrite, gr3
 234 => b"00010_0010_01_000000000000", -- add, gr2
 235 => b"00000_0000_00_000000000001", -- 1
 236 => b"10000_0010_00_000000000000", -- tpoint, gr2
 237 => b"01111_0000_00_000000000000", -- tread, gr0
 238 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 239 => b"00110_0000_01_000000000000", -- beq
 240 => b"00000_0000_00_000011111010", -- P1LEFT
 241 => b"01110_0011_00_000000000000", -- twrite, gr3
 242 => b"00010_0010_01_000000000000", -- add, gr2
 243 => b"00000_0000_00_000000000001", -- 1
 244 => b"10000_0010_00_000000000000", -- tpoint, gr2
 245 => b"01111_0000_00_000000000000", -- tread, gr0
 246 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 247 => b"00110_0000_01_000000000000", -- beq
 248 => b"00000_0000_00_000011111010", -- P1LEFT
 249 => b"01110_0011_00_000000000000", -- twrite, gr3
 250 => b"00000_0010_00_001011101100", -- load, gr2, P1BOMB1POS
 251 => b"00011_0010_01_000000000000", -- sub, gr2
 252 => b"00000_0000_00_000000000001", -- 1
 253 => b"10000_0010_00_000000000000", -- tpoint, gr2
 254 => b"01111_0000_00_000000000000", -- tread, gr0
 255 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 256 => b"00110_0000_01_000000000000", -- beq
 257 => b"00000_0000_00_000100001011", -- P1DOWN
 258 => b"01110_0011_00_000000000000", -- twrite, gr3
 259 => b"00011_0010_01_000000000000", -- sub, gr2
 260 => b"00000_0000_00_000000000001", -- 1
 261 => b"10000_0010_00_000000000000", -- tpoint, gr2
 262 => b"01111_0000_00_000000000000", -- tread, gr0
 263 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 264 => b"00110_0000_01_000000000000", -- beq
 265 => b"00000_0000_00_000100001011", -- P1DOWN
 266 => b"01110_0011_00_000000000000", -- twrite, gr3
 267 => b"00000_0010_00_001011101100", -- load, gr2, P1BOMB1POS
 268 => b"00010_0010_01_000000000000", -- add, gr2
 269 => b"00000_0000_00_000000001111", -- 15
 270 => b"10000_0010_00_000000000000", -- tpoint, gr2
 271 => b"01111_0000_00_000000000000", -- tread, gr0
 272 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 273 => b"00110_0000_01_000000000000", -- beq
 274 => b"00000_0000_00_000100011100", -- P1UP
 275 => b"01110_0011_00_000000000000", -- twrite, gr3
 276 => b"00010_0010_01_000000000000", -- add, gr2
 277 => b"00000_0000_00_000000001111", -- 15
 278 => b"10000_0010_00_000000000000", -- tpoint, gr2
 279 => b"01111_0000_00_000000000000", -- tread, gr0
 280 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 281 => b"00110_0000_01_000000000000", -- beq
 282 => b"00000_0000_00_000100011100", -- P1UP
 283 => b"01110_0011_00_000000000000", -- twrite, gr3
 284 => b"00000_0010_00_001011101100", -- load, gr2, P1BOMB1POS
 285 => b"00011_0010_01_000000000000", -- sub, gr2
 286 => b"00000_0000_00_000000001111", -- 15
 287 => b"10000_0010_00_000000000000", -- tpoint, gr2
 288 => b"01111_0000_00_000000000000", -- tread, gr0
 289 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 290 => b"00110_0000_01_000000000000", -- beq
 291 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 292 => b"01110_0011_00_000000000000", -- twrite, gr3
 293 => b"00011_0010_01_000000000000", -- sub, gr2
 294 => b"00000_0000_00_000000001111", -- 15
 295 => b"10000_0010_00_000000000000", -- tpoint, gr2
 296 => b"01111_0000_00_000000000000", -- tread, gr0
 297 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 298 => b"00110_0000_01_000000000000", -- beq
 299 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 300 => b"01110_0011_00_000000000000", -- twrite, gr3
 301 => b"00100_0000_01_000000000000", -- jump
 302 => b"00000_0000_00_000011000110", -- TICKBOMB1_R
 303 => b"00000_0000_00_001100000000", -- load, gr0, P2BOMB1ACTIVE
 304 => b"00011_0000_01_000000000000", -- sub, gr0
 305 => b"00000_0000_00_000000000001", -- 1
 306 => b"00111_0000_01_000000000000", -- bne
 307 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 308 => b"00000_0000_00_001011111111", -- load, gr0, P2BOMB1TIME
 309 => b"00011_0000_01_000000000000", -- sub, gr0
 310 => b"00000_0000_00_000000000001", -- 1
 311 => b"00001_0000_10_001011111111", -- store, gr0, P2BOMB1TIME
 312 => b"00000_0000_01_000000000000", -- load, gr0
 313 => b"00000_0000_00_000000000000", -- 0
 314 => b"00011_0000_00_001011111111", -- sub, gr0, P2BOMB1TIME
 315 => b"00110_0000_01_000000000000", -- beq
 316 => b"00000_0000_00_000100111111", -- EXPLODE2
 317 => b"00100_0000_01_000000000000", -- jump
 318 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 319 => b"00000_0000_00_001011111110", -- load, gr0, P2BOMB1POS
 320 => b"00001_0000_10_001100000011", -- store, gr0, P2EXPLOSION1POS
 321 => b"00000_0000_01_000000000000", -- load, gr0
 322 => b"00000_0000_00_000000000001", -- 1
 323 => b"00001_0000_10_001100000010", -- store, gr0, P2EXPLOSION1ACTIVE
 324 => b"00000_0000_01_000000000000", -- load, gr0
 325 => b"00000_0000_00_000000000010", -- 2
 326 => b"00001_0000_10_001100000001", -- store, gr0, P2EXPLOSION1TIME
 327 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 328 => b"00011_0000_01_000000000000", -- sub, gr0
 329 => b"00000_0000_00_000000000001", -- 1
 330 => b"00001_0000_10_001100010001", -- store, gr0, P2BOMBCOUNT
 331 => b"00000_0010_00_001011111110", -- load, gr2, P2BOMB1POS
 332 => b"00000_0011_00_001100011101", -- load, gr3, EXPLOSION
 333 => b"10000_0010_00_000000000000", -- tpoint, gr2
 334 => b"01110_0011_00_000000000000", -- twrite, gr3
 335 => b"00010_0010_01_000000000000", -- add, gr2
 336 => b"00000_0000_00_000000000001", -- 1
 337 => b"10000_0010_00_000000000000", -- tpoint, gr2
 338 => b"01111_0000_00_000000000000", -- tread, gr0
 339 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 340 => b"00110_0000_01_000000000000", -- beq
 341 => b"00000_0000_00_000101011111", -- P2LEFT
 342 => b"01110_0011_00_000000000000", -- twrite, gr3
 343 => b"00010_0010_01_000000000000", -- add, gr2
 344 => b"00000_0000_00_000000000001", -- 1
 345 => b"10000_0010_00_000000000000", -- tpoint, gr2
 346 => b"01111_0000_00_000000000000", -- tread, gr0
 347 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 348 => b"00110_0000_01_000000000000", -- beq
 349 => b"00000_0000_00_000101011111", -- P2LEFT
 350 => b"01110_0011_00_000000000000", -- twrite, gr3
 351 => b"00000_0010_00_001011111110", -- load, gr2, P2BOMB1POS
 352 => b"00011_0010_01_000000000000", -- sub, gr2
 353 => b"00000_0000_00_000000000001", -- 1
 354 => b"10000_0010_00_000000000000", -- tpoint, gr2
 355 => b"01111_0000_00_000000000000", -- tread, gr0
 356 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 357 => b"00110_0000_01_000000000000", -- beq
 358 => b"00000_0000_00_000101110000", -- P2DOWN
 359 => b"01110_0011_00_000000000000", -- twrite, gr3
 360 => b"00011_0010_01_000000000000", -- sub, gr2
 361 => b"00000_0000_00_000000000001", -- 1
 362 => b"10000_0010_00_000000000000", -- tpoint, gr2
 363 => b"01111_0000_00_000000000000", -- tread, gr0
 364 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 365 => b"00110_0000_01_000000000000", -- beq
 366 => b"00000_0000_00_000101110000", -- P2DOWN
 367 => b"01110_0011_00_000000000000", -- twrite, gr3
 368 => b"00000_0010_00_001011111110", -- load, gr2, P2BOMB1POS
 369 => b"00010_0010_01_000000000000", -- add, gr2
 370 => b"00000_0000_00_000000001111", -- 15
 371 => b"10000_0010_00_000000000000", -- tpoint, gr2
 372 => b"01111_0000_00_000000000000", -- tread, gr0
 373 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 374 => b"00110_0000_01_000000000000", -- beq
 375 => b"00000_0000_00_000110000001", -- P2UP
 376 => b"01110_0011_00_000000000000", -- twrite, gr3
 377 => b"00010_0010_01_000000000000", -- add, gr2
 378 => b"00000_0000_00_000000001111", -- 15
 379 => b"10000_0010_00_000000000000", -- tpoint, gr2
 380 => b"01111_0000_00_000000000000", -- tread, gr0
 381 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 382 => b"00110_0000_01_000000000000", -- beq
 383 => b"00000_0000_00_000110000001", -- P2UP
 384 => b"01110_0011_00_000000000000", -- twrite, gr3
 385 => b"00000_0010_00_001011111110", -- load, gr2, P2BOMB1POS
 386 => b"00011_0010_01_000000000000", -- sub, gr2
 387 => b"00000_0000_00_000000001111", -- 15
 388 => b"10000_0010_00_000000000000", -- tpoint, gr2
 389 => b"01111_0000_00_000000000000", -- tread, gr0
 390 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 391 => b"00110_0000_01_000000000000", -- beq
 392 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 393 => b"01110_0011_00_000000000000", -- twrite, gr3
 394 => b"00011_0010_01_000000000000", -- sub, gr2
 395 => b"00000_0000_00_000000001111", -- 15
 396 => b"10000_0010_00_000000000000", -- tpoint, gr2
 397 => b"01111_0000_00_000000000000", -- tread, gr0
 398 => b"00011_0000_00_001100011011", -- sub, gr0, WALL
 399 => b"00110_0000_01_000000000000", -- beq
 400 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 401 => b"01110_0011_00_000000000000", -- twrite, gr3
 402 => b"00100_0000_01_000000000000", -- jump
 403 => b"00000_0000_00_000011001000", -- TICKBOMB2_R
 404 => b"10101_0000_01_000000000000", -- btn1
 405 => b"00000_0000_00_000110011010", -- BTN1
 406 => b"11010_0000_01_000000000000", -- btn2
 407 => b"00000_0000_00_000111110100", -- BTN2
 408 => b"00100_0000_01_000000000000", -- jump
 409 => b"00000_0000_00_000000000100", -- BUTTON_R
 410 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 411 => b"00011_0000_00_001100010010", -- sub, gr0, MAXBOMBS
 412 => b"00110_0000_01_000000000000", -- beq
 413 => b"00000_0000_00_000110010110", -- BTN1_R
 414 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 415 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 416 => b"00000_0000_00_001100010100", -- load, gr0, YPOS1
 417 => b"01000_0000_01_000000000000", -- mul, gr0
 418 => b"00000_0000_00_000000001111", -- 15
 419 => b"00010_0000_00_001100010011", -- add, gr0, XPOS1
 420 => b"10000_0000_00_000000000000", -- tpoint, gr0
 421 => b"01111_0001_00_000000000000", -- tread, gr1
 422 => b"00011_0001_00_001100011110", -- sub, gr1, EGG
 423 => b"00110_0000_01_000000000000", -- beq
 424 => b"00000_0000_00_000110010110", -- BTN1_R
 425 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 426 => b"00011_0000_01_000000000000", -- sub, gr0
 427 => b"00000_0000_00_000000000000", -- 0
 428 => b"00110_0000_01_000000000000", -- beq
 429 => b"00000_0000_00_000110111110", -- P1PLACEBOMB1
 430 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 431 => b"00011_0000_01_000000000000", -- sub, gr0
 432 => b"00000_0000_00_000000000001", -- 1
 433 => b"00110_0000_01_000000000000", -- beq
 434 => b"00000_0000_00_000111010000", -- P1PLACEBOMB2
 435 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 436 => b"00011_0000_01_000000000000", -- sub, gr0
 437 => b"00000_0000_00_000000000010", -- 2
 438 => b"00110_0000_01_000000000000", -- beq
 439 => b"00000_0000_00_000111010000", -- P1PLACEBOMB2
 440 => b"00000_0000_00_001100010000", -- load, gr0, P1BOMBCOUNT
 441 => b"00010_0000_01_000000000000", -- add, gr0
 442 => b"00000_0000_00_000000000001", -- 1
 443 => b"00001_0000_10_001100010000", -- store, gr0, P1BOMBCOUNT
 444 => b"00100_0000_01_000000000000", -- jump
 445 => b"00000_0000_00_000110010110", -- BTN1_R
 446 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 447 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 448 => b"00000_0011_00_001100010100", -- load, gr3, YPOS1
 449 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 450 => b"01000_0011_01_000000000000", -- mul, gr3
 451 => b"00000_0000_00_000000001111", -- 15
 452 => b"00010_0011_00_001100010011", -- add, gr3, XPOS1
 453 => b"10000_0011_00_000000000000", -- tpoint, gr3
 454 => b"01110_0010_00_000000000000", -- twrite, gr2
 455 => b"00000_0000_01_000000000000", -- load, gr0
 456 => b"00000_0000_00_000000000001", -- 1
 457 => b"00001_0000_10_001011101110", -- store, gr0, P1BOMB1ACTIVE
 458 => b"00001_0011_10_001011101100", -- store, gr3, P1BOMB1POS
 459 => b"00000_0000_01_000000000000", -- load, gr0
 460 => b"00000_0000_00_000000010000", -- 16
 461 => b"00001_0000_10_001011101101", -- store, gr0, P1BOMB1TIME
 462 => b"00100_0000_01_000000000000", -- jump
 463 => b"00000_0000_00_000110111000", -- P1INCREASEBOMBCOUNTER
 464 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 465 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 466 => b"00000_0011_00_001100010100", -- load, gr3, YPOS1
 467 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 468 => b"01000_0011_01_000000000000", -- mul, gr3
 469 => b"00000_0000_00_000000001111", -- 15
 470 => b"00010_0011_00_001100010011", -- add, gr3, XPOS1
 471 => b"10000_0011_00_000000000000", -- tpoint, gr3
 472 => b"01110_0010_00_000000000000", -- twrite, gr2
 473 => b"00000_0000_01_000000000000", -- load, gr0
 474 => b"00000_0000_00_000000000001", -- 1
 475 => b"00001_0000_10_001011110100", -- store, gr0, P1BOMB2ACTIVE
 476 => b"00001_0011_10_001011110010", -- store, gr3, P1BOMB2POS
 477 => b"00000_0000_01_000000000000", -- load, gr0
 478 => b"00000_0000_00_000000010000", -- 16
 479 => b"00001_0000_10_001011110011", -- store, gr0, P1BOMB2TIME
 480 => b"00100_0000_01_000000000000", -- jump
 481 => b"00000_0000_00_000110111000", -- P1INCREASEBOMBCOUNTER
 482 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 483 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 484 => b"00000_0011_00_001100010100", -- load, gr3, YPOS1
 485 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 486 => b"01000_0011_01_000000000000", -- mul, gr3
 487 => b"00000_0000_00_000000001111", -- 15
 488 => b"00010_0011_00_001100010011", -- add, gr3, XPOS1
 489 => b"10000_0011_00_000000000000", -- tpoint, gr3
 490 => b"01110_0010_00_000000000000", -- twrite, gr2
 491 => b"00000_0000_01_000000000000", -- load, gr0
 492 => b"00000_0000_00_000000000001", -- 1
 493 => b"00001_0000_10_001011111010", -- store, gr0, P1BOMB3ACTIVE
 494 => b"00001_0011_10_001011111000", -- store, gr3, P1BOMB3POS
 495 => b"00000_0000_01_000000000000", -- load, gr0
 496 => b"00000_0000_00_000000010000", -- 16
 497 => b"00001_0000_10_001011111001", -- store, gr0, P1BOMB3TIME
 498 => b"00100_0000_01_000000000000", -- jump
 499 => b"00000_0000_00_000110111000", -- P1INCREASEBOMBCOUNTER
 500 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 501 => b"00011_0000_00_001100010010", -- sub, gr0, MAXBOMBS
 502 => b"00110_0000_01_000000000000", -- beq
 503 => b"00000_0000_00_000110011000", -- BTN2_R
 504 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 505 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 506 => b"00000_0000_00_001100010110", -- load, gr0, YPOS2
 507 => b"01000_0000_01_000000000000", -- mul, gr0
 508 => b"00000_0000_00_000000001111", -- 15
 509 => b"00010_0000_00_001100010101", -- add, gr0, XPOS2
 510 => b"10000_0000_00_000000000000", -- tpoint, gr0
 511 => b"01111_0001_00_000000000000", -- tread, gr1
 512 => b"00011_0001_00_001100011110", -- sub, gr1, EGG
 513 => b"00110_0000_01_000000000000", -- beq
 514 => b"00000_0000_00_000110011000", -- BTN2_R
 515 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 516 => b"00011_0000_01_000000000000", -- sub, gr0
 517 => b"00000_0000_00_000000000000", -- 0
 518 => b"00110_0000_01_000000000000", -- beq
 519 => b"00000_0000_00_001000011000", -- P2PLACEBOMB1
 520 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 521 => b"00011_0000_01_000000000000", -- sub, gr0
 522 => b"00000_0000_00_000000000001", -- 1
 523 => b"00110_0000_01_000000000000", -- beq
 524 => b"00000_0000_00_001000101010", -- P2PLACEBOMB2
 525 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 526 => b"00011_0000_01_000000000000", -- sub, gr0
 527 => b"00000_0000_00_000000000010", -- 2
 528 => b"00110_0000_01_000000000000", -- beq
 529 => b"00000_0000_00_001000111100", -- P2PLACEBOMB3
 530 => b"00000_0000_00_001100010001", -- load, gr0, P2BOMBCOUNT
 531 => b"00010_0000_01_000000000000", -- add, gr0
 532 => b"00000_0000_00_000000000001", -- 1
 533 => b"00001_0000_10_001100010001", -- store, gr0, P2BOMBCOUNT
 534 => b"00100_0000_01_000000000000", -- jump
 535 => b"00000_0000_00_000110011000", -- BTN2_R
 536 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 537 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 538 => b"00000_0011_00_001100010110", -- load, gr3, YPOS2
 539 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 540 => b"01000_0011_01_000000000000", -- mul, gr3
 541 => b"00000_0000_00_000000001111", -- 15
 542 => b"00010_0011_00_001100010101", -- add, gr3, XPOS2
 543 => b"10000_0011_00_000000000000", -- tpoint, gr3
 544 => b"01110_0010_00_000000000000", -- twrite, gr2
 545 => b"00000_0000_01_000000000000", -- load, gr0
 546 => b"00000_0000_00_000000000001", -- 1
 547 => b"00001_0000_10_001100000000", -- store, gr0, P2BOMB1ACTIVE
 548 => b"00001_0011_10_001011111110", -- store, gr3, P2BOMB1POS
 549 => b"00000_0000_01_000000000000", -- load, gr0
 550 => b"00000_0000_00_000000010000", -- 16
 551 => b"00001_0000_10_001011111111", -- store, gr0, P2BOMB1TIME
 552 => b"00100_0000_01_000000000000", -- jump
 553 => b"00000_0000_00_001000010010", -- P2INCREASEBOMBCOUNTER
 554 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 555 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 556 => b"00000_0011_00_001100010110", -- load, gr3, YPOS2
 557 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 558 => b"01000_0011_01_000000000000", -- mul, gr3
 559 => b"00000_0000_00_000000001111", -- 15
 560 => b"00010_0011_00_001100010101", -- add, gr3, XPOS2
 561 => b"10000_0011_00_000000000000", -- tpoint, gr3
 562 => b"01110_0010_00_000000000000", -- twrite, gr2
 563 => b"00000_0000_01_000000000000", -- load, gr0
 564 => b"00000_0000_00_000000000001", -- 1
 565 => b"00001_0000_10_001100000110", -- store, gr0, P2BOMB2ACTIVE
 566 => b"00001_0011_10_001100000100", -- store, gr3, P2BOMB2POS
 567 => b"00000_0000_01_000000000000", -- load, gr0
 568 => b"00000_0000_00_000000010000", -- 16
 569 => b"00001_0000_10_001100000101", -- store, gr0, P2BOMB2TIME
 570 => b"00100_0000_01_000000000000", -- jump
 571 => b"00000_0000_00_001000010010", -- P2INCREASEBOMBCOUNTER
 572 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 573 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 574 => b"00000_0011_00_001100010110", -- load, gr3, YPOS2
 575 => b"00000_0010_00_001100011110", -- load, gr2, EGG
 576 => b"01000_0011_01_000000000000", -- mul, gr3
 577 => b"00000_0000_00_000000001111", -- 15
 578 => b"00010_0011_00_001100010101", -- add, gr3, XPOS2
 579 => b"10000_0011_00_000000000000", -- tpoint, gr3
 580 => b"01110_0010_00_000000000000", -- twrite, gr2
 581 => b"00000_0000_01_000000000000", -- load, gr0
 582 => b"00000_0000_00_000000000001", -- 1
 583 => b"00001_0000_10_001100001100", -- store, gr0, P2BOMB3ACTIVE
 584 => b"00001_0011_10_001100001010", -- store, gr3, P2BOMB3POS
 585 => b"00000_0000_01_000000000000", -- load, gr0
 586 => b"00000_0000_00_000000010000", -- 16
 587 => b"00001_0000_10_001100001011", -- store, gr0, P2BOMB3TIME
 588 => b"00100_0000_01_000000000000", -- jump
 589 => b"00000_0000_00_001000010010", -- P2INCREASEBOMBCOUNTER
 590 => b"00100_0000_01_000000000000", -- jump
 591 => b"00000_0000_00_001011101010", -- COUNT1
 592 => b"10001_0000_01_000000000000", -- joy1r
 593 => b"00000_0000_00_001001100010", -- P1R
 594 => b"10011_0000_01_000000000000", -- joy1l
 595 => b"00000_0000_00_001010000100", -- P1L
 596 => b"10010_0000_01_000000000000", -- joy1u
 597 => b"00000_0000_00_001001110011", -- P1U
 598 => b"10100_0000_01_000000000000", -- joy1d
 599 => b"00000_0000_00_001010010101", -- P1D
 600 => b"10110_0000_01_000000000000", -- joy2r
 601 => b"00000_0000_00_001010100110", -- P2R
 602 => b"11000_0000_01_000000000000", -- joy2l
 603 => b"00000_0000_00_001011001000", -- P2L
 604 => b"10111_0000_01_000000000000", -- joy2u
 605 => b"00000_0000_00_001010110111", -- P2U
 606 => b"11001_0000_01_000000000000", -- joy2d
 607 => b"00000_0000_00_001011011001", -- P2D
 608 => b"00100_0000_01_000000000000", -- jump
 609 => b"00000_0000_00_000000000010", -- CONTROL_R
 610 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 611 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 612 => b"00000_0000_00_001100010100", -- load, gr0, YPOS1
 613 => b"01000_0000_01_000000000000", -- mul, gr0
 614 => b"00000_0000_00_000000001111", -- 15
 615 => b"00010_0000_00_001100010011", -- add, gr0, XPOS1
 616 => b"00010_0000_01_000000000000", -- add, gr0
 617 => b"00000_0000_00_000000000001", -- 1
 618 => b"10000_0000_00_000000000000", -- tpoint, gr0
 619 => b"01111_0001_00_000000000000", -- tread, gr1
 620 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 621 => b"00111_0000_01_000000000000", -- bne
 622 => b"00000_0000_00_001001010100", -- J1
 623 => b"00010_1100_01_000000000000", -- add, gr12
 624 => b"00000_0000_00_000000000001", -- 1
 625 => b"00100_0000_01_000000000000", -- jump
 626 => b"00000_0000_00_001001010100", -- J1
 627 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 628 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 629 => b"00000_0000_00_001100010100", -- load, gr0, YPOS1
 630 => b"00011_0000_01_000000000000", -- sub, gr0
 631 => b"00000_0000_00_000000000001", -- 1
 632 => b"01000_0000_01_000000000000", -- mul, gr0
 633 => b"00000_0000_00_000000001111", -- 15
 634 => b"00010_0000_00_001100010011", -- add, gr0, XPOS1
 635 => b"10000_0000_00_000000000000", -- tpoint, gr0
 636 => b"01111_0001_00_000000000000", -- tread, gr1
 637 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 638 => b"00111_0000_01_000000000000", -- bne
 639 => b"00000_0000_00_001001011000", -- J2
 640 => b"00011_1101_01_000000000000", -- sub, gr13
 641 => b"00000_0000_00_000000000001", -- 1
 642 => b"00100_0000_01_000000000000", -- jump
 643 => b"00000_0000_00_001001011000", -- J2
 644 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 645 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 646 => b"00000_0000_00_001100010100", -- load, gr0, YPOS1
 647 => b"01000_0000_01_000000000000", -- mul, gr0
 648 => b"00000_0000_00_000000001111", -- 15
 649 => b"00010_0000_00_001100010011", -- add, gr0, XPOS1
 650 => b"00011_0000_01_000000000000", -- sub, gr0
 651 => b"00000_0000_00_000000000001", -- 1
 652 => b"10000_0000_00_000000000000", -- tpoint, gr0
 653 => b"01111_0001_00_000000000000", -- tread, gr1
 654 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 655 => b"00111_0000_01_000000000000", -- bne
 656 => b"00000_0000_00_001001010100", -- J1
 657 => b"00011_1100_01_000000000000", -- sub, gr12
 658 => b"00000_0000_00_000000000001", -- 1
 659 => b"00100_0000_01_000000000000", -- jump
 660 => b"00000_0000_00_001001010100", -- J1
 661 => b"00001_1100_10_001100010011", -- store, gr12, XPOS1
 662 => b"00001_1101_10_001100010100", -- store, gr13, YPOS1
 663 => b"00000_0000_00_001100010100", -- load, gr0, YPOS1
 664 => b"00010_0000_01_000000000000", -- add, gr0
 665 => b"00000_0000_00_000000000001", -- 1
 666 => b"01000_0000_01_000000000000", -- mul, gr0
 667 => b"00000_0000_00_000000001111", -- 15
 668 => b"00010_0000_00_001100010011", -- add, gr0, XPOS1
 669 => b"10000_0000_00_000000000000", -- tpoint, gr0
 670 => b"01111_0001_00_000000000000", -- tread, gr1
 671 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 672 => b"00111_0000_01_000000000000", -- bne
 673 => b"00000_0000_00_001001011000", -- J2
 674 => b"00010_1101_01_000000000000", -- add, gr13
 675 => b"00000_0000_00_000000000001", -- 1
 676 => b"00100_0000_01_000000000000", -- jump
 677 => b"00000_0000_00_001001011000", -- J2
 678 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 679 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 680 => b"00000_0000_00_001100010110", -- load, gr0, YPOS2
 681 => b"01000_0000_01_000000000000", -- mul, gr0
 682 => b"00000_0000_00_000000001111", -- 15
 683 => b"00010_0000_00_001100010101", -- add, gr0, XPOS2
 684 => b"00010_0000_01_000000000000", -- add, gr0
 685 => b"00000_0000_00_000000000001", -- 1
 686 => b"10000_0000_00_000000000000", -- tpoint, gr0
 687 => b"01111_0001_00_000000000000", -- tread, gr1
 688 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 689 => b"00111_0000_01_000000000000", -- bne
 690 => b"00000_0000_00_001001011100", -- J3
 691 => b"00010_1110_01_000000000000", -- add, gr14
 692 => b"00000_0000_00_000000000001", -- 1
 693 => b"00100_0000_01_000000000000", -- jump
 694 => b"00000_0000_00_001001011100", -- J3
 695 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 696 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 697 => b"00000_0000_00_001100010110", -- load, gr0, YPOS2
 698 => b"00011_0000_01_000000000000", -- sub, gr0
 699 => b"00000_0000_00_000000000001", -- 1
 700 => b"01000_0000_01_000000000000", -- mul, gr0
 701 => b"00000_0000_00_000000001111", -- 15
 702 => b"00010_0000_00_001100010101", -- add, gr0, XPOS2
 703 => b"10000_0000_00_000000000000", -- tpoint, gr0
 704 => b"01111_0001_00_000000000000", -- tread, gr1
 705 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 706 => b"00111_0000_01_000000000000", -- bne
 707 => b"00000_0000_00_000000000010", -- CONTROL_R
 708 => b"00011_1111_01_000000000000", -- sub, gr15
 709 => b"00000_0000_00_000000000001", -- 1
 710 => b"00100_0000_01_000000000000", -- jump
 711 => b"00000_0000_00_000000000010", -- CONTROL_R
 712 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 713 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 714 => b"00000_0000_00_001100010110", -- load, gr0, YPOS2
 715 => b"01000_0000_01_000000000000", -- mul, gr0
 716 => b"00000_0000_00_000000001111", -- 15
 717 => b"00010_0000_00_001100010101", -- add, gr0, XPOS2
 718 => b"00011_0000_01_000000000000", -- sub, gr0
 719 => b"00000_0000_00_000000000001", -- 1
 720 => b"10000_0000_00_000000000000", -- tpoint, gr0
 721 => b"01111_0001_00_000000000000", -- tread, gr1
 722 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 723 => b"00111_0000_01_000000000000", -- bne
 724 => b"00000_0000_00_001001011100", -- J3
 725 => b"00011_1110_01_000000000000", -- sub, gr14
 726 => b"00000_0000_00_000000000001", -- 1
 727 => b"00100_0000_01_000000000000", -- jump
 728 => b"00000_0000_00_001001011100", -- J3
 729 => b"00001_1110_10_001100010101", -- store, gr14, XPOS2
 730 => b"00001_1111_10_001100010110", -- store, gr15, YPOS2
 731 => b"00000_0000_00_001100010110", -- load, gr0, YPOS2
 732 => b"00010_0000_01_000000000000", -- add, gr0
 733 => b"00000_0000_00_000000000001", -- 1
 734 => b"01000_0000_01_000000000000", -- mul, gr0
 735 => b"00000_0000_00_000000001111", -- 15
 736 => b"00010_0000_00_001100010101", -- add, gr0, XPOS2
 737 => b"10000_0000_00_000000000000", -- tpoint, gr0
 738 => b"01111_0001_00_000000000000", -- tread, gr1
 739 => b"00011_0001_00_001100011010", -- sub, gr1, GRASS
 740 => b"00111_0000_01_000000000000", -- bne
 741 => b"00000_0000_00_000000000010", -- CONTROL_R
 742 => b"00010_1111_01_000000000000", -- add, gr15
 743 => b"00000_0000_00_000000000001", -- 1
 744 => b"00100_0000_01_000000000000", -- jump
 745 => b"00000_0000_00_000000000010", -- CONTROL_R
 746 => b"00100_0000_01_000000000000", -- jump
 747 => b"00000_0000_00_001001010000", -- COUNT_R
 748 => b"00000_0000_00_000000000000", -- 0
 749 => b"00000_0000_00_000000000000", -- 0
 750 => b"00000_0000_00_000000000000", -- 0
 751 => b"00000_0000_00_000000000000", -- 0
 752 => b"00000_0000_00_000000000000", -- 0
 753 => b"00000_0000_00_000000000000", -- 0
 754 => b"00000_0000_00_000000000000", -- 0
 755 => b"00000_0000_00_000000000000", -- 0
 756 => b"00000_0000_00_000000000000", -- 0
 757 => b"00000_0000_00_000000000000", -- 0
 758 => b"00000_0000_00_000000000000", -- 0
 759 => b"00000_0000_00_000000000000", -- 0
 760 => b"00000_0000_00_000000000000", -- 0
 761 => b"00000_0000_00_000000000000", -- 0
 762 => b"00000_0000_00_000000000000", -- 0
 763 => b"00000_0000_00_000000000000", -- 0
 764 => b"00000_0000_00_000000000000", -- 0
 765 => b"00000_0000_00_000000000000", -- 0
 766 => b"00000_0000_00_000000000000", -- 0
 767 => b"00000_0000_00_000000000000", -- 0
 768 => b"00000_0000_00_000000000000", -- 0
 769 => b"00000_0000_00_000000000000", -- 0
 770 => b"00000_0000_00_000000000000", -- 0
 771 => b"00000_0000_00_000000000000", -- 0
 772 => b"00000_0000_00_000000000000", -- 0
 773 => b"00000_0000_00_000000000000", -- 0
 774 => b"00000_0000_00_000000000000", -- 0
 775 => b"00000_0000_00_000000000000", -- 0
 776 => b"00000_0000_00_000000000000", -- 0
 777 => b"00000_0000_00_000000000000", -- 0
 778 => b"00000_0000_00_000000000000", -- 0
 779 => b"00000_0000_00_000000000000", -- 0
 780 => b"00000_0000_00_000000000000", -- 0
 781 => b"00000_0000_00_000000000000", -- 0
 782 => b"00000_0000_00_000000000000", -- 0
 783 => b"00000_0000_00_000000000000", -- 0
 784 => b"00000_0000_00_000000000000", -- 0
 785 => b"00000_0000_00_000000000000", -- 0
 786 => b"00000_0000_00_000000000011", -- 3
 787 => b"00000_0000_00_000000000000", -- 0
 788 => b"00000_0000_00_000000000000", -- 0
 789 => b"00000_0000_00_000000000000", -- 0
 790 => b"00000_0000_00_000000000000", -- 0
 791 => b"00000_0000_00_000000000000", -- 0
 792 => b"00000_0000_00_000000000000", -- 0
 793 => b"00000_0000_00_000000000000", -- 0
 794 => b"00000_0000_00_000000000000", -- 0
 795 => b"00000_0000_00_000000000001", -- 1
 796 => b"00000_0000_00_000000000010", -- 2
 797 => b"00000_0000_00_000000000011", -- 3
 798 => b"00000_0000_00_000000000100", -- 4


    others => (others => '0')
  );

  signal PM : pm_t := pm_c;


begin  -- pMem

  PM_out <= PM(to_integer(pAddr));

  process (clk)
  begin
    if rising_edge(clk) then
      if PM_write = '1' then
        PM(to_integer(pAddr)) <= PM_in;
      end if;
    end if;
  end process;
  
 -- PM(to_integer(pAddr)) <= PM_in when PM_write = '1' else PM(to_integer(pAddr));

end Behavioral; 
